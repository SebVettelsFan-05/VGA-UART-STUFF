module image_rom (
	input logic [9:0] v_count,
	input logic [9:0] h_count,
	output logic [11:0] rgb_colour
);
	logic [9:0] v_count_n;
	logic [9:0] h_count_n;
	assign v_count_n = v_count >> 2;
	assign h_count_n = h_count >> 2;

	logic [11:0] array[0:19199] = '{
		12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h344, 12'h444, 12'h334, 12'h444, 12'h444, 12'h334, 12'h344, 12'h444, 12'h434, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h455, 12'h455, 12'h445, 12'h444, 12'h455, 12'h545, 12'h455, 12'h555, 12'h555, 12'h454, 12'h555, 12'h555, 12'h455, 12'h555, 12'h545, 12'h455, 12'h555, 12'h545, 12'h444, 12'h555, 12'h545, 12'h444, 12'h545, 12'h544, 12'h444, 12'h555, 12'h444, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h566, 12'h556, 12'h566, 12'h565, 12'h556, 12'h665, 12'h566, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h445, 12'h455, 12'h554, 12'h444, 12'h555, 12'h445, 12'h544, 12'h555, 12'h444, 12'h444, 12'h544, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h545, 12'h444, 12'h544, 12'h444, 12'h444, 12'h445,
		12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h434, 12'h344, 12'h444, 12'h433, 12'h334, 12'h444, 12'h333, 12'h333, 12'h444, 12'h444, 12'h334, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h455, 12'h444, 12'h454, 12'h555, 12'h444, 12'h554, 12'h455, 12'h544, 12'h444, 12'h445, 12'h555, 12'h444, 12'h555, 12'h545, 12'h445, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h455, 12'h554, 12'h454, 12'h445, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h565, 12'h555, 12'h666, 12'h665, 12'h556, 12'h556, 12'h565, 12'h666, 12'h566, 12'h565, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h554, 12'h445, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h444, 12'h555, 12'h545, 12'h445, 12'h554, 12'h545, 12'h545, 12'h455, 12'h555, 12'h544, 12'h555, 12'h455, 12'h545, 12'h555, 12'h444, 12'h544, 12'h545, 12'h454, 12'h455,
		12'h444, 12'h454, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h344, 12'h445, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h443, 12'h434, 12'h433, 12'h343, 12'h444, 12'h434, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h455, 12'h444, 12'h454, 12'h455, 12'h445, 12'h554, 12'h455, 12'h545, 12'h455, 12'h554, 12'h545, 12'h454, 12'h555, 12'h545, 12'h454, 12'h555, 12'h555, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h554, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h554, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h565, 12'h565, 12'h556, 12'h566, 12'h556, 12'h565, 12'h656, 12'h566, 12'h565, 12'h656, 12'h566, 12'h556, 12'h655, 12'h666, 12'h566, 12'h566, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h566, 12'h556, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h445, 12'h555, 12'h555, 12'h445, 12'h545, 12'h555, 12'h444, 12'h555, 12'h555, 12'h444, 12'h555, 12'h454, 12'h544, 12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h444, 12'h454, 12'h555, 12'h544, 12'h455, 12'h555, 12'h555,
		12'h445, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h334, 12'h344, 12'h444, 12'h434, 12'h344, 12'h444, 12'h434, 12'h344, 12'h444, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h455, 12'h444, 12'h445, 12'h455, 12'h545, 12'h455, 12'h555, 12'h455, 12'h455, 12'h445, 12'h454, 12'h555, 12'h445, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h545, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h455, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h555, 12'h565, 12'h566, 12'h666, 12'h555, 12'h566, 12'h666, 12'h666, 12'h565, 12'h666, 12'h566, 12'h555, 12'h655, 12'h566, 12'h556, 12'h565, 12'h566, 12'h666, 12'h555, 12'h565, 12'h556, 12'h555, 12'h565, 12'h556, 12'h555, 12'h566, 12'h555, 12'h566, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h544, 12'h555, 12'h455, 12'h544, 12'h555, 12'h455, 12'h545, 12'h454, 12'h555, 12'h444, 12'h554, 12'h455, 12'h544, 12'h555, 12'h555, 12'h544, 12'h445, 12'h554, 12'h445, 12'h544, 12'h555, 12'h555,
		12'h445, 12'h454, 12'h445, 12'h445, 12'h444, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h334, 12'h344, 12'h444, 12'h444, 12'h444, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h445, 12'h445, 12'h444, 12'h445, 12'h454, 12'h444, 12'h445, 12'h454, 12'h444, 12'h455, 12'h445, 12'h454, 12'h455, 12'h445, 12'h554, 12'h555, 12'h455, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h454, 12'h545, 12'h455, 12'h454, 12'h545, 12'h445, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h444, 12'h444, 12'h444, 12'h434, 12'h444, 12'h444, 12'h444, 12'h334, 12'h444, 12'h444, 12'h333, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h545, 12'h555, 12'h444, 12'h445, 12'h555, 12'h555, 12'h555, 12'h566, 12'h566, 12'h656, 12'h565, 12'h556, 12'h665, 12'h566, 12'h656, 12'h556, 12'h666, 12'h666, 12'h566, 12'h555, 12'h666, 12'h656, 12'h566, 12'h566, 12'h656, 12'h566, 12'h566, 12'h656, 12'h555, 12'h566, 12'h555, 12'h555, 12'h565, 12'h555, 12'h556, 12'h566, 12'h555, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h544, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h554, 12'h555, 12'h555, 12'h555, 12'h454, 12'h445, 12'h555, 12'h555, 12'h555,
		12'h454, 12'h455, 12'h444, 12'h455, 12'h445, 12'h454, 12'h455, 12'h455, 12'h445, 12'h455, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h433, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h445, 12'h454, 12'h455, 12'h445, 12'h444, 12'h455, 12'h444, 12'h455, 12'h445, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h434, 12'h434, 12'h344, 12'h333, 12'h333, 12'h334, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h434, 12'h433, 12'h333, 12'h334, 12'h434, 12'h333, 12'h333, 12'h444, 12'h434, 12'h433, 12'h444, 12'h334, 12'h455, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h556, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h556, 12'h565, 12'h565, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h665, 12'h656, 12'h566, 12'h555, 12'h566, 12'h556, 12'h565, 12'h565, 12'h556, 12'h565, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555,
		12'h445, 12'h455, 12'h444, 12'h445, 12'h455, 12'h444, 12'h444, 12'h444, 12'h455, 12'h455, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h434, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h455, 12'h554, 12'h554, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h454, 12'h445, 12'h444, 12'h454, 12'h445, 12'h545, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h455, 12'h555, 12'h445, 12'h455, 12'h544, 12'h545, 12'h444, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h444, 12'h434, 12'h333, 12'h444, 12'h433, 12'h333, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h434, 12'h444, 12'h444, 12'h333, 12'h444, 12'h444, 12'h555, 12'h565, 12'h666, 12'h555, 12'h666, 12'h666, 12'h665, 12'h666, 12'h566, 12'h666, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h566, 12'h656, 12'h666, 12'h565, 12'h556, 12'h566, 12'h556, 12'h555, 12'h566, 12'h556, 12'h555, 12'h566, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h554, 12'h545, 12'h555, 12'h444, 12'h555,
		12'h455, 12'h555, 12'h455, 12'h445, 12'h445, 12'h455, 12'h444, 12'h445, 12'h455, 12'h444, 12'h444, 12'h454, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h554, 12'h455, 12'h445, 12'h555, 12'h445, 12'h554, 12'h555, 12'h444, 12'h554, 12'h555, 12'h445, 12'h455, 12'h555, 12'h454, 12'h454, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h434, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h222, 12'h222, 12'h323, 12'h222, 12'h323, 12'h333, 12'h333, 12'h333, 12'h222, 12'h333, 12'h333, 12'h333, 12'h323, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h333, 12'h332, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h545, 12'h555, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h565, 12'h555, 12'h566, 12'h555, 12'h566, 12'h565, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h455, 12'h555, 12'h554, 12'h455, 12'h455, 12'h555, 12'h455, 12'h444, 12'h445, 12'h455, 12'h445, 12'h454, 12'h454, 12'h445, 12'h454, 12'h445, 12'h445, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h445, 12'h455, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h223, 12'h223, 12'h222, 12'h333, 12'h223, 12'h222, 12'h333, 12'h222, 12'h333, 12'h322, 12'h222, 12'h333, 12'h333, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h323, 12'h222, 12'h333, 12'h222, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h444, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h665, 12'h666, 12'h556, 12'h655, 12'h665, 12'h665, 12'h566, 12'h666, 12'h555, 12'h556, 12'h655, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h445, 12'h455, 12'h455, 12'h445, 12'h454, 12'h455, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h454, 12'h445, 12'h445, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h566, 12'h555, 12'h555, 12'h444, 12'h334, 12'h434, 12'h344, 12'h544, 12'h444, 12'h333, 12'h434, 12'h333, 12'h434, 12'h433, 12'h323, 12'h333, 12'h222, 12'h332, 12'h333, 12'h333, 12'h333, 12'h323, 12'h444, 12'h333, 12'h322, 12'h222, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h222, 12'h333, 12'h333, 12'h222, 12'h222, 12'h333, 12'h222, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h444, 12'h445, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h656, 12'h566, 12'h655, 12'h656, 12'h565, 12'h666, 12'h666, 12'h656, 12'h556, 12'h556, 12'h655, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h455, 12'h555, 12'h455, 12'h445, 12'h555, 12'h455, 12'h444, 12'h555, 12'h455, 12'h554, 12'h555, 12'h445, 12'h555, 12'h455, 12'h445, 12'h455, 12'h454, 12'h455, 12'h445, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h455, 12'h544, 12'h445, 12'h555, 12'h454, 12'h555, 12'h555, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h444, 12'h344, 12'h333, 12'h444, 12'h333, 12'h333, 12'h333, 12'h434, 12'h333, 12'h444, 12'h333, 12'h333, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h333, 12'h332, 12'h222, 12'h222, 12'h222, 12'h223, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h323, 12'h333, 12'h223, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h333, 12'h323, 12'h333, 12'h333, 12'h333, 12'h222, 12'h333, 12'h333, 12'h343, 12'h555, 12'h445, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h565, 12'h566, 12'h666, 12'h666, 12'h566, 12'h566, 12'h666, 12'h555, 12'h656, 12'h666, 12'h665, 12'h566, 12'h666, 12'h666, 12'h566, 12'h656, 12'h656, 12'h656, 12'h555, 12'h666, 12'h656, 12'h566, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h455, 12'h445, 12'h455, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h455, 12'h445, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h322, 12'h333, 12'h332, 12'h323, 12'h333, 12'h333, 12'h323, 12'h322, 12'h222, 12'h333, 12'h222, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h323, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h333, 12'h333, 12'h443, 12'h455, 12'h555, 12'h666, 12'h666, 12'h677, 12'h676, 12'h666, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h566, 12'h566, 12'h665, 12'h566, 12'h666, 12'h655, 12'h566, 12'h665, 12'h656, 12'h666, 12'h555, 12'h555, 12'h555, 12'h566, 12'h566, 12'h666, 12'h566, 12'h566, 12'h666, 12'h555, 12'h555,
		12'h455, 12'h445, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h455, 12'h555, 12'h555, 12'h555, 12'h545, 12'h454, 12'h455, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h566, 12'h566, 12'h566, 12'h666, 12'h566, 12'h555, 12'h445, 12'h444, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h322, 12'h433, 12'h333, 12'h333, 12'h322, 12'h333, 12'h434, 12'h333, 12'h333, 12'h333, 12'h322, 12'h332, 12'h322, 12'h323, 12'h333, 12'h333, 12'h222, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h323, 12'h222, 12'h222, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h222, 12'h222, 12'h233, 12'h333, 12'h555, 12'h666, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h665, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h556, 12'h555, 12'h666, 12'h565, 12'h656, 12'h656, 12'h655, 12'h555, 12'h665, 12'h655, 12'h566, 12'h666, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h455, 12'h555, 12'h455, 12'h555, 12'h455, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h444, 12'h454, 12'h555, 12'h545, 12'h445, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h555, 12'h566, 12'h566, 12'h565, 12'h555, 12'h545, 12'h444, 12'h334, 12'h444, 12'h434, 12'h333, 12'h444, 12'h434, 12'h333, 12'h333, 12'h333, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h333, 12'h333, 12'h322, 12'h222, 12'h332, 12'h222, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h222, 12'h222, 12'h222, 12'h121, 12'h222, 12'h222, 12'h112, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h444, 12'h444, 12'h666, 12'h666, 12'h766, 12'h777, 12'h677, 12'h666, 12'h677, 12'h666, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h656, 12'h565, 12'h566, 12'h555, 12'h656, 12'h556, 12'h565, 12'h656, 12'h555, 12'h666, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h566, 12'h565, 12'h566, 12'h566, 12'h566, 12'h565, 12'h656, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h333, 12'h444, 12'h444, 12'h333, 12'h333, 12'h434, 12'h444, 12'h333, 12'h433, 12'h323, 12'h333, 12'h444, 12'h444, 12'h433, 12'h333, 12'h333, 12'h433, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h322, 12'h333, 12'h333, 12'h333, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h111, 12'h212, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h444, 12'h666, 12'h666, 12'h666, 12'h776, 12'h777, 12'h666, 12'h666, 12'h677, 12'h667, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h656, 12'h666, 12'h655, 12'h566, 12'h666, 12'h656, 12'h566, 12'h666, 12'h565, 12'h656, 12'h565, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h455, 12'h455, 12'h555, 12'h455, 12'h455, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h666, 12'h566, 12'h566, 12'h655, 12'h555, 12'h445, 12'h444, 12'h444, 12'h434, 12'h444, 12'h333, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h434, 12'h444, 12'h444, 12'h434, 12'h333, 12'h433, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h444, 12'h544, 12'h544, 12'h443, 12'h544, 12'h544, 12'h543, 12'h543, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h121, 12'h111, 12'h111, 12'h211, 12'h111, 12'h111, 12'h211, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h333, 12'h555, 12'h666, 12'h666, 12'h777, 12'h666, 12'h677, 12'h666, 12'h777, 12'h676, 12'h676, 12'h677, 12'h666, 12'h677, 12'h677, 12'h666, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h656, 12'h666, 12'h665, 12'h555, 12'h656, 12'h666, 12'h555, 12'h566, 12'h666, 12'h555, 12'h566,
		12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h566, 12'h566, 12'h556, 12'h666, 12'h666, 12'h566, 12'h665, 12'h666, 12'h656, 12'h666, 12'h666, 12'h566, 12'h555, 12'h544, 12'h444, 12'h344, 12'h334, 12'h444, 12'h333, 12'h223, 12'h222, 12'h223, 12'h322, 12'h333, 12'h444, 12'h434, 12'h444, 12'h544, 12'h555, 12'h444, 12'h544, 12'h544, 12'h544, 12'h544, 12'h434, 12'h433, 12'h433, 12'h543, 12'h544, 12'h544, 12'h544, 12'h654, 12'h644, 12'h644, 12'h544, 12'h544, 12'h543, 12'h533, 12'h533, 12'h533, 12'h644, 12'h533, 12'h433, 12'h432, 12'h433, 12'h432, 12'h422, 12'h432, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h221, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h211, 12'h111, 12'h111, 12'h221, 12'h211, 12'h222, 12'h111, 12'h222, 12'h444, 12'h555, 12'h666, 12'h677, 12'h676, 12'h777, 12'h767, 12'h666, 12'h766, 12'h776, 12'h776, 12'h667, 12'h766, 12'h676, 12'h777, 12'h667, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666,
		12'h555, 12'h455, 12'h555, 12'h556, 12'h556, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h455, 12'h556, 12'h555, 12'h455, 12'h556, 12'h555, 12'h455, 12'h555, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h566, 12'h556, 12'h565, 12'h666, 12'h656, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h555, 12'h666, 12'h545, 12'h555, 12'h444, 12'h444, 12'h444, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h222, 12'h323, 12'h333, 12'h333, 12'h433, 12'h545, 12'h544, 12'h544, 12'h544, 12'h544, 12'h544, 12'h654, 12'h544, 12'h544, 12'h544, 12'h544, 12'h433, 12'h544, 12'h544, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h643, 12'h644, 12'h644, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h433, 12'h332, 12'h433, 12'h322, 12'h322, 12'h322, 12'h222, 12'h322, 12'h222, 12'h222, 12'h211, 12'h121, 12'h222, 12'h211, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h212, 12'h221, 12'h222, 12'h111, 12'h222, 12'h222, 12'h112, 12'h122, 12'h221, 12'h222, 12'h222, 12'h222, 12'h666, 12'h666, 12'h777, 12'h777, 12'h677, 12'h777, 12'h677, 12'h767, 12'h667, 12'h666, 12'h766, 12'h666, 12'h767, 12'h776, 12'h666, 12'h677, 12'h676, 12'h666, 12'h677, 12'h676, 12'h666, 12'h666, 12'h676, 12'h666, 12'h666, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h666, 12'h656, 12'h665, 12'h566, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666,
		12'h555, 12'h555, 12'h556, 12'h565, 12'h556, 12'h556, 12'h555, 12'h556, 12'h455, 12'h555, 12'h456, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h556, 12'h566, 12'h566, 12'h565, 12'h556, 12'h666, 12'h666, 12'h566, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h555, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h434, 12'h433, 12'h434, 12'h333, 12'h333, 12'h322, 12'h222, 12'h233, 12'h333, 12'h222, 12'h333, 12'h433, 12'h444, 12'h544, 12'h555, 12'h655, 12'h755, 12'h765, 12'h755, 12'h755, 12'h654, 12'h755, 12'h644, 12'h655, 12'h644, 12'h654, 12'h644, 12'h755, 12'h755, 12'h754, 12'h754, 12'h754, 12'h744, 12'h754, 12'h643, 12'h744, 12'h744, 12'h744, 12'h643, 12'h643, 12'h743, 12'h743, 12'h643, 12'h743, 12'h643, 12'h533, 12'h543, 12'h533, 12'h433, 12'h432, 12'h432, 12'h433, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h211, 12'h221, 12'h211, 12'h221, 12'h222, 12'h222, 12'h221, 12'h111, 12'h111, 12'h122, 12'h212, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h111, 12'h111, 12'h111, 12'h333, 12'h555, 12'h666, 12'h777, 12'h677, 12'h777, 12'h676, 12'h777, 12'h677, 12'h777, 12'h677, 12'h666, 12'h777, 12'h666, 12'h666, 12'h767, 12'h677, 12'h766, 12'h677, 12'h777, 12'h666, 12'h777, 12'h677, 12'h676, 12'h676, 12'h676, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666,
		12'h556, 12'h556, 12'h566, 12'h565, 12'h556, 12'h565, 12'h565, 12'h556, 12'h455, 12'h555, 12'h555, 12'h456, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h566, 12'h556, 12'h555, 12'h566, 12'h555, 12'h566, 12'h566, 12'h566, 12'h565, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h556, 12'h444, 12'h445, 12'h444, 12'h444, 12'h555, 12'h555, 12'h444, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h222, 12'h434, 12'h433, 12'h333, 12'h434, 12'h544, 12'h544, 12'h655, 12'h766, 12'h877, 12'h877, 12'h866, 12'h976, 12'h855, 12'h855, 12'h754, 12'h754, 12'h755, 12'h855, 12'h865, 12'h855, 12'h754, 12'h754, 12'h754, 12'h854, 12'h854, 12'h854, 12'h854, 12'h754, 12'h743, 12'h854, 12'h753, 12'h743, 12'h744, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h643, 12'h633, 12'h633, 12'h543, 12'h533, 12'h433, 12'h432, 12'h532, 12'h432, 12'h432, 12'h432, 12'h422, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h111, 12'h222, 12'h222, 12'h221, 12'h111, 12'h222, 12'h222, 12'h211, 12'h121, 12'h211, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h444, 12'h666, 12'h776, 12'h666, 12'h777, 12'h776, 12'h776, 12'h777, 12'h777, 12'h776, 12'h777, 12'h777, 12'h776, 12'h777, 12'h666, 12'h666, 12'h777, 12'h666, 12'h777, 12'h677, 12'h766, 12'h777, 12'h677, 12'h777, 12'h777, 12'h676, 12'h676, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676,
		12'h555, 12'h566, 12'h566, 12'h556, 12'h566, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h455, 12'h556, 12'h556, 12'h565, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h666, 12'h566, 12'h666, 12'h656, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h555, 12'h444, 12'h444, 12'h444, 12'h434, 12'h434, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h434, 12'h444, 12'h655, 12'h766, 12'h866, 12'h877, 12'h988, 12'hA88, 12'h977, 12'hA77, 12'h976, 12'h976, 12'h976, 12'h965, 12'h865, 12'h966, 12'h965, 12'h965, 12'h965, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h955, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h753, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h632, 12'h643, 12'h633, 12'h633, 12'h543, 12'h633, 12'h533, 12'h533, 12'h532, 12'h432, 12'h432, 12'h432, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h211, 12'h211, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h444, 12'h555, 12'h666, 12'h666, 12'h667, 12'h777, 12'h777, 12'h667, 12'h776, 12'h767, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676,
		12'h565, 12'h566, 12'h555, 12'h566, 12'h566, 12'h556, 12'h566, 12'h566, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h566, 12'h556, 12'h566, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h556, 12'h655, 12'h545, 12'h555, 12'h445, 12'h333, 12'h444, 12'h333, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h655, 12'h766, 12'h877, 12'hA98, 12'hA88, 12'hB99, 12'hA99, 12'hA88, 12'hA88, 12'hA87, 12'hA88, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h965, 12'h965, 12'h954, 12'h954, 12'h954, 12'h954, 12'h964, 12'h954, 12'h965, 12'h954, 12'h954, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h844, 12'h844, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h532, 12'h533, 12'h533, 12'h532, 12'h432, 12'h432, 12'h432, 12'h422, 12'h322, 12'h322, 12'h322, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h122, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h223, 12'h334, 12'h666, 12'h666, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h767, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676, 12'h676,
		12'h556, 12'h556, 12'h566, 12'h566, 12'h556, 12'h565, 12'h566, 12'h556, 12'h565, 12'h566, 12'h556, 12'h566, 12'h555, 12'h566, 12'h566, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h677, 12'h677, 12'h667, 12'h676, 12'h777, 12'h555, 12'h444, 12'h444, 12'h545, 12'h545, 12'h444, 12'h333, 12'h333, 12'h334, 12'h333, 12'h333, 12'h334, 12'h333, 12'h333, 12'h434, 12'h434, 12'h554, 12'h766, 12'h988, 12'hA99, 12'hB99, 12'hBAA, 12'hBAA, 12'hC99, 12'hCAA, 12'hBA9, 12'hB99, 12'hB88, 12'hB88, 12'hA87, 12'hA77, 12'hB87, 12'hA87, 12'hA76, 12'hA76, 12'h976, 12'hA65, 12'h965, 12'h965, 12'h965, 12'h965, 12'h965, 12'h964, 12'h964, 12'h965, 12'h954, 12'h954, 12'h954, 12'h854, 12'h854, 12'h854, 12'h743, 12'h753, 12'h743, 12'h743, 12'h643, 12'h743, 12'h643, 12'h643, 12'h743, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h533, 12'h532, 12'h532, 12'h433, 12'h432, 12'h432, 12'h432, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h211, 12'h222, 12'h111, 12'h222, 12'h112, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h344, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h676, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h766, 12'h666, 12'h666, 12'h666, 12'h676, 12'h676, 12'h676, 12'h777, 12'h777,
		12'h556, 12'h565, 12'h566, 12'h556, 12'h665, 12'h566, 12'h556, 12'h556, 12'h565, 12'h556, 12'h566, 12'h566, 12'h555, 12'h556, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h676, 12'h667, 12'h677, 12'h677, 12'h677, 12'h666, 12'h666, 12'h555, 12'h556, 12'h555, 12'h555, 12'h544, 12'h444, 12'h333, 12'h333, 12'h333, 12'h334, 12'h444, 12'h333, 12'h433, 12'h434, 12'h444, 12'h444, 12'h867, 12'hA99, 12'hBAA, 12'hBAA, 12'hCBB, 12'hCCC, 12'hCBB, 12'hCBA, 12'hCBB, 12'hB99, 12'hC99, 12'hCAA, 12'hB98, 12'hB88, 12'hB88, 12'hB98, 12'hB87, 12'hB87, 12'hA76, 12'hA76, 12'hA76, 12'hA65, 12'hA65, 12'hA65, 12'hA76, 12'hA65, 12'h965, 12'h954, 12'h964, 12'h954, 12'h954, 12'h954, 12'h954, 12'h954, 12'h854, 12'h854, 12'h854, 12'h743, 12'h744, 12'h743, 12'h743, 12'h643, 12'h633, 12'h643, 12'h643, 12'h643, 12'h633, 12'h633, 12'h532, 12'h533, 12'h533, 12'h532, 12'h532, 12'h433, 12'h432, 12'h433, 12'h432, 12'h432, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h221, 12'h222, 12'h111, 12'h111, 12'h211, 12'h222, 12'h222, 12'h221, 12'h112, 12'h222, 12'h111, 12'h111, 12'h222, 12'h555, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h777, 12'h787, 12'h787, 12'h777, 12'h787, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h677, 12'h777, 12'h776, 12'h777, 12'h767, 12'h777, 12'h776, 12'h777, 12'h777,
		12'h556, 12'h565, 12'h556, 12'h656, 12'h566, 12'h656, 12'h566, 12'h565, 12'h556, 12'h555, 12'h566, 12'h556, 12'h566, 12'h565, 12'h556, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h677, 12'h676, 12'h677, 12'h667, 12'h676, 12'h677, 12'h667, 12'h777, 12'h777, 12'h666, 12'h666, 12'h555, 12'h444, 12'h545, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h334, 12'h444, 12'h433, 12'h333, 12'h444, 12'h434, 12'h544, 12'h644, 12'h655, 12'hA88, 12'hBAA, 12'hCBB, 12'hCBB, 12'hDBB, 12'hDCC, 12'hDBB, 12'hCBB, 12'hDBB, 12'hDBB, 12'hDBA, 12'hCA9, 12'hB98, 12'hC98, 12'hB87, 12'hC99, 12'hB88, 12'hB87, 12'hB76, 12'hA76, 12'hA75, 12'hA75, 12'hA65, 12'hA75, 12'hA65, 12'hA76, 12'hA65, 12'h965, 12'h965, 12'h955, 12'h965, 12'h964, 12'h954, 12'h954, 12'h854, 12'h854, 12'h844, 12'h853, 12'h743, 12'h744, 12'h744, 12'h643, 12'h744, 12'h743, 12'h743, 12'h643, 12'h643, 12'h643, 12'h533, 12'h532, 12'h533, 12'h533, 12'h533, 12'h532, 12'h432, 12'h433, 12'h432, 12'h432, 12'h432, 12'h432, 12'h322, 12'h322, 12'h332, 12'h322, 12'h222, 12'h221, 12'h122, 12'h221, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h211, 12'h111, 12'h111, 12'h222, 12'h566, 12'h777, 12'h777, 12'h777, 12'h787, 12'h777, 12'h777, 12'h787, 12'h777, 12'h777, 12'h787, 12'h787, 12'h787, 12'h787, 12'h777, 12'h788, 12'h887, 12'h888, 12'h787, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h676, 12'h666, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777,
		12'h566, 12'h556, 12'h665, 12'h566, 12'h556, 12'h565, 12'h656, 12'h566, 12'h556, 12'h566, 12'h555, 12'h555, 12'h566, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h677, 12'h666, 12'h777, 12'h676, 12'h666, 12'h555, 12'h555, 12'h444, 12'h434, 12'h555, 12'h666, 12'h444, 12'h434, 12'h434, 12'h333, 12'h444, 12'h545, 12'h434, 12'h333, 12'h444, 12'h433, 12'h544, 12'h655, 12'h977, 12'hBAA, 12'hCBB, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDBB, 12'hDCC, 12'hCBB, 12'hCAA, 12'hB99, 12'hB98, 12'hC98, 12'hC98, 12'hB87, 12'hB87, 12'hB86, 12'hB76, 12'hA65, 12'hA66, 12'hA76, 12'hA76, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'hA65, 12'h954, 12'h965, 12'h964, 12'h954, 12'h954, 12'h954, 12'h854, 12'h854, 12'h843, 12'h743, 12'h744, 12'h743, 12'h744, 12'h743, 12'h633, 12'h643, 12'h643, 12'h643, 12'h533, 12'h532, 12'h532, 12'h533, 12'h532, 12'h533, 12'h533, 12'h532, 12'h433, 12'h433, 12'h432, 12'h432, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h222, 12'h211, 12'h121, 12'h111, 12'h112, 12'h121, 12'h211, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h444, 12'h665, 12'h676, 12'h777, 12'h787, 12'h888, 12'h888, 12'h788, 12'h888, 12'h788, 12'h778, 12'h787, 12'h878, 12'h778, 12'h887, 12'h877, 12'h778, 12'h888, 12'h878, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h677, 12'h776, 12'h777, 12'h777, 12'h777,
		12'h566, 12'h656, 12'h566, 12'h566, 12'h556, 12'h565, 12'h556, 12'h556, 12'h665, 12'h556, 12'h566, 12'h666, 12'h656, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h677, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h556, 12'h555, 12'h545, 12'h444, 12'h444, 12'h555, 12'h656, 12'h544, 12'h444, 12'h444, 12'h333, 12'h444, 12'h555, 12'h444, 12'h333, 12'h433, 12'h444, 12'h554, 12'h755, 12'h877, 12'hBAA, 12'hBAA, 12'hCBC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDBB, 12'hDBB, 12'hDBB, 12'hDCB, 12'hDBB, 12'hDBA, 12'hC99, 12'hC99, 12'hB87, 12'hB87, 12'hB87, 12'hB77, 12'hB87, 12'hB76, 12'hA76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA75, 12'hA76, 12'hA65, 12'hA65, 12'hA65, 12'h954, 12'h964, 12'h955, 12'hA65, 12'h954, 12'h965, 12'h954, 12'h954, 12'h954, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h532, 12'h533, 12'h532, 12'h533, 12'h532, 12'h432, 12'h423, 12'h432, 12'h432, 12'h422, 12'h432, 12'h332, 12'h322, 12'h322, 12'h322, 12'h222, 12'h221, 12'h221, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h444, 12'h677, 12'h777, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h877, 12'h788, 12'h777, 12'h888, 12'h888, 12'h787, 12'h887, 12'h888, 12'h788, 12'h887, 12'h777, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h677, 12'h777, 12'h777,
		12'h566, 12'h656, 12'h565, 12'h556, 12'h666, 12'h666, 12'h566, 12'h565, 12'h656, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676, 12'h677, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h666, 12'h545, 12'h445, 12'h666, 12'h444, 12'h555, 12'h555, 12'h555, 12'h444, 12'h434, 12'h333, 12'h434, 12'h555, 12'h444, 12'h333, 12'h434, 12'h444, 12'h434, 12'h655, 12'h877, 12'hBAA, 12'hCBB, 12'hDBC, 12'hDCC, 12'hCBB, 12'hCBA, 12'hCAA, 12'hDBB, 12'hCAA, 12'hDBA, 12'hDAA, 12'hCAA, 12'hCA9, 12'hC98, 12'hB87, 12'hC88, 12'hB87, 12'hB87, 12'hB76, 12'hB87, 12'hB76, 12'hB87, 12'hB76, 12'hB76, 12'hB76, 12'hB75, 12'hB75, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'hA64, 12'hA65, 12'hA65, 12'h964, 12'h954, 12'h965, 12'h964, 12'h954, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h743, 12'h743, 12'h633, 12'h633, 12'h643, 12'h532, 12'h533, 12'h543, 12'h533, 12'h532, 12'h533, 12'h532, 12'h432, 12'h433, 12'h433, 12'h432, 12'h433, 12'h433, 12'h332, 12'h333, 12'h322, 12'h322, 12'h222, 12'h222, 12'h221, 12'h111, 12'h222, 12'h211, 12'h222, 12'h222, 12'h111, 12'h221, 12'h222, 12'h222, 12'h444, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h887, 12'h777, 12'h887, 12'h778, 12'h778, 12'h887, 12'h777, 12'h788, 12'h877, 12'h787, 12'h788, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h566, 12'h566, 12'h656, 12'h565, 12'h666, 12'h556, 12'h565, 12'h566, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h667, 12'h677, 12'h677, 12'h777, 12'h777, 12'h677, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h666, 12'h777, 12'h555, 12'h555, 12'h666, 12'h555, 12'h545, 12'h555, 12'h666, 12'h545, 12'h444, 12'h545, 12'h444, 12'h666, 12'h545, 12'h433, 12'h444, 12'h433, 12'h444, 12'h544, 12'h877, 12'hA88, 12'hB99, 12'hCBB, 12'hDBA, 12'hDAA, 12'hCAA, 12'hDBA, 12'hDBB, 12'hCBA, 12'hDAA, 12'hDAA, 12'hCA9, 12'hC99, 12'hC88, 12'hC98, 12'hC87, 12'hC98, 12'hB87, 12'hC87, 12'hB76, 12'hC87, 12'hB77, 12'hB75, 12'hB75, 12'hB76, 12'hA65, 12'hB76, 12'hB75, 12'hA65, 12'hA65, 12'hA65, 12'h955, 12'hA65, 12'hA65, 12'h954, 12'h965, 12'h955, 12'h965, 12'h965, 12'h954, 12'h954, 12'h854, 12'h854, 12'h854, 12'h844, 12'h744, 12'h744, 12'h744, 12'h743, 12'h643, 12'h643, 12'h532, 12'h533, 12'h532, 12'h532, 12'h643, 12'h533, 12'h533, 12'h532, 12'h432, 12'h422, 12'h422, 12'h432, 12'h433, 12'h422, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h211, 12'h222, 12'h122, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h444, 12'h666, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h887, 12'h888, 12'h878, 12'h887, 12'h778, 12'h887, 12'h878, 12'h777, 12'h887, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h556, 12'h666, 12'h566, 12'h656, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h667, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h677, 12'h666, 12'h555, 12'h544, 12'h444, 12'h656, 12'h655, 12'h545, 12'h445, 12'h545, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h444, 12'h656, 12'h544, 12'h444, 12'h433, 12'h533, 12'h544, 12'h866, 12'hA88, 12'hCA9, 12'hCAA, 12'hCAA, 12'hDAA, 12'hDA9, 12'hDBA, 12'hDBB, 12'hCAA, 12'hDBA, 12'hDAA, 12'hCA9, 12'hC98, 12'hC88, 12'hC98, 12'hC88, 12'hB76, 12'hC87, 12'hB76, 12'hC87, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'h965, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'h955, 12'h954, 12'h854, 12'h854, 12'h955, 12'h854, 12'h854, 12'h753, 12'h744, 12'h754, 12'h743, 12'h643, 12'h643, 12'h633, 12'h643, 12'h643, 12'h532, 12'h533, 12'h533, 12'h532, 12'h532, 12'h432, 12'h433, 12'h432, 12'h322, 12'h432, 12'h432, 12'h433, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h122, 12'h222, 12'h111, 12'h111, 12'h212, 12'h344, 12'h666, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h887, 12'h778, 12'h887, 12'h787, 12'h878, 12'h787, 12'h877, 12'h878, 12'h788, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h566, 12'h656, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h777, 12'h788, 12'h777, 12'h555, 12'h545, 12'h444, 12'h444, 12'h445, 12'h545, 12'h444, 12'h555, 12'h434, 12'h545, 12'h555, 12'h555, 12'h444, 12'h434, 12'h444, 12'h555, 12'h444, 12'h544, 12'h544, 12'h544, 12'h755, 12'h865, 12'hA77, 12'hB87, 12'hC98, 12'hC99, 12'hCA9, 12'hDAA, 12'hC99, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC99, 12'hCA9, 12'hC98, 12'hC98, 12'hB87, 12'hB76, 12'hB76, 12'hC87, 12'hB76, 12'hC76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hC76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA75, 12'hA65, 12'hB65, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'h954, 12'h964, 12'h965, 12'h854, 12'h854, 12'h853, 12'h854, 12'h744, 12'h643, 12'h643, 12'h643, 12'h633, 12'h643, 12'h533, 12'h643, 12'h532, 12'h533, 12'h532, 12'h432, 12'h433, 12'h432, 12'h422, 12'h433, 12'h322, 12'h322, 12'h433, 12'h332, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h444, 12'h666, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h878, 12'h878, 12'h888, 12'h877, 12'h878, 12'h887, 12'h877, 12'h788, 12'h787, 12'h777, 12'h878, 12'h787, 12'h877, 12'h888, 12'h787, 12'h787, 12'h777, 12'h787, 12'h787, 12'h777, 12'h777,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h788, 12'h888, 12'h888, 12'h888, 12'h666, 12'h555, 12'h545, 12'h444, 12'h545, 12'h555, 12'h555, 12'h555, 12'h444, 12'h666, 12'h777, 12'h655, 12'h555, 12'h544, 12'h333, 12'h555, 12'h655, 12'h655, 12'h655, 12'h544, 12'h644, 12'h644, 12'h866, 12'h976, 12'hB87, 12'hC98, 12'hC98, 12'hDBA, 12'hDAA, 12'hDA9, 12'hDBA, 12'hDBA, 12'hCAA, 12'hDAA, 12'hDA9, 12'hD98, 12'hC88, 12'hC87, 12'hB76, 12'hC87, 12'hC87, 12'hC76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC86, 12'hC76, 12'hB76, 12'hC76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'hB76, 12'hB75, 12'hA65, 12'hA65, 12'hB75, 12'hB75, 12'hA65, 12'h955, 12'h964, 12'h965, 12'h965, 12'h954, 12'h854, 12'h854, 12'h843, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h633, 12'h633, 12'h642, 12'h633, 12'h533, 12'h533, 12'h532, 12'h422, 12'h422, 12'h432, 12'h433, 12'h432, 12'h422, 12'h322, 12'h333, 12'h322, 12'h332, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h121, 12'h111, 12'h222, 12'h666, 12'h888, 12'h888, 12'h898, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h877, 12'h878, 12'h887, 12'h878, 12'h787, 12'h788, 12'h877, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h777,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h676, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h788, 12'h788, 12'h888, 12'h888, 12'h777, 12'h555, 12'h555, 12'h444, 12'h444, 12'h555, 12'h545, 12'h555, 12'h655, 12'h767, 12'h555, 12'h777, 12'h656, 12'h655, 12'h544, 12'h434, 12'h555, 12'h656, 12'h655, 12'h544, 12'h555, 12'h655, 12'h755, 12'h866, 12'h977, 12'hB88, 12'hB99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDBA, 12'hDA9, 12'hC99, 12'hC98, 12'hC88, 12'hC87, 12'hC87, 12'hC87, 12'hB77, 12'hC76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC86, 12'hC86, 12'hB76, 12'hB76, 12'hA66, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'h965, 12'h954, 12'h955, 12'h964, 12'h954, 12'h954, 12'h854, 12'h854, 12'h743, 12'h744, 12'h743, 12'h643, 12'h633, 12'h643, 12'h532, 12'h633, 12'h532, 12'h533, 12'h532, 12'h532, 12'h532, 12'h432, 12'h432, 12'h433, 12'h432, 12'h432, 12'h433, 12'h322, 12'h332, 12'h323, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h112, 12'h555, 12'h777, 12'h888, 12'h888, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h877, 12'h877, 12'h788, 12'h877, 12'h888, 12'h788, 12'h877, 12'h788, 12'h877, 12'h777, 12'h888, 12'h888, 12'h787, 12'h777,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h788, 12'h788, 12'h887, 12'h888, 12'h788, 12'h788, 12'h777, 12'h655, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h555, 12'h656, 12'h777, 12'h777, 12'h766, 12'h655, 12'h656, 12'h555, 12'h545, 12'h444, 12'h656, 12'h544, 12'h544, 12'h655, 12'h655, 12'h755, 12'h865, 12'hA76, 12'hB87, 12'hC98, 12'hC98, 12'hDA9, 12'hDBA, 12'hDAA, 12'hDAA, 12'hD99, 12'hDA9, 12'hD99, 12'hC97, 12'hC87, 12'hC88, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA76, 12'hB76, 12'hB75, 12'hB76, 12'hA76, 12'hA65, 12'hA65, 12'h954, 12'h965, 12'h955, 12'h954, 12'h854, 12'h854, 12'h744, 12'h744, 12'h743, 12'h643, 12'h633, 12'h643, 12'h643, 12'h632, 12'h643, 12'h643, 12'h632, 12'h533, 12'h532, 12'h533, 12'h432, 12'h422, 12'h422, 12'h422, 12'h433, 12'h432, 12'h422, 12'h433, 12'h333, 12'h322, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h222, 12'h666, 12'h777, 12'h888, 12'h998, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h787, 12'h878, 12'h888, 12'h888, 12'h888, 12'h887, 12'h777, 12'h788, 12'h787, 12'h777, 12'h888, 12'h788,
		12'h666, 12'h667, 12'h667, 12'h667, 12'h666, 12'h667, 12'h667, 12'h666, 12'h667, 12'h766, 12'h766, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h788, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h555, 12'h666, 12'h555, 12'h445, 12'h555, 12'h878, 12'h767, 12'h666, 12'h766, 12'h767, 12'h656, 12'h544, 12'h555, 12'h545, 12'h544, 12'h544, 12'h555, 12'h655, 12'h544, 12'h655, 12'h644, 12'h755, 12'h855, 12'hA77, 12'hB87, 12'hC88, 12'hC98, 12'hDA9, 12'hDAA, 12'hDBA, 12'hDA9, 12'hD98, 12'hC98, 12'hC98, 12'hD98, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC77, 12'hC87, 12'hD87, 12'hD97, 12'hD97, 12'hD97, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hB76, 12'hC87, 12'hB86, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'hA65, 12'h964, 12'h965, 12'h955, 12'h954, 12'h854, 12'h854, 12'h744, 12'h743, 12'h743, 12'h643, 12'h643, 12'h633, 12'h533, 12'h533, 12'h532, 12'h533, 12'h533, 12'h532, 12'h533, 12'h432, 12'h432, 12'h433, 12'h432, 12'h422, 12'h332, 12'h432, 12'h322, 12'h332, 12'h333, 12'h332, 12'h322, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h222, 12'h343, 12'h777, 12'h888, 12'h888, 12'h888, 12'h999, 12'h998, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h877, 12'h778, 12'h788, 12'h888,
		12'h666, 12'h666, 12'h677, 12'h776, 12'h677, 12'h667, 12'h777, 12'h777, 12'h667, 12'h777, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h666, 12'h545, 12'h555, 12'h556, 12'h767, 12'h777, 12'h878, 12'h878, 12'h776, 12'h767, 12'h655, 12'h766, 12'h555, 12'h555, 12'h544, 12'h544, 12'h544, 12'h544, 12'h544, 12'h756, 12'h644, 12'h654, 12'h654, 12'h855, 12'hA66, 12'hB87, 12'hB88, 12'hC98, 12'hC98, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA8, 12'hD98, 12'hD98, 12'hD98, 12'hC97, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC76, 12'hC86, 12'hC76, 12'hC86, 12'hC86, 12'hC76, 12'hB76, 12'hB75, 12'hA65, 12'hA65, 12'h965, 12'hA65, 12'h965, 12'h965, 12'h954, 12'h854, 12'h754, 12'h743, 12'h743, 12'h743, 12'h743, 12'h643, 12'h633, 12'h643, 12'h633, 12'h532, 12'h532, 12'h532, 12'h533, 12'h532, 12'h533, 12'h533, 12'h432, 12'h432, 12'h423, 12'h332, 12'h432, 12'h433, 12'h322, 12'h322, 12'h322, 12'h232, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h111, 12'h111, 12'h121, 12'h222, 12'h333, 12'h777, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h888, 12'h888, 12'h888, 12'h887, 12'h878, 12'h778, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h787, 12'h788, 12'h777, 12'h787,
		12'h767, 12'h777, 12'h766, 12'h767, 12'h777, 12'h766, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h666, 12'h556, 12'h656, 12'h656, 12'h777, 12'h555, 12'h777, 12'h777, 12'h988, 12'h655, 12'h666, 12'h666, 12'h666, 12'h767, 12'h655, 12'h655, 12'h554, 12'h644, 12'h655, 12'h654, 12'h755, 12'h755, 12'h866, 12'h865, 12'h965, 12'hA76, 12'hB76, 12'hC87, 12'hC88, 12'hC98, 12'hD98, 12'hD98, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD87, 12'hD87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hB87, 12'hB87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC77, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC86, 12'hC87, 12'hB76, 12'hA75, 12'hA65, 12'h964, 12'hA65, 12'h965, 12'h965, 12'h954, 12'h854, 12'h854, 12'h743, 12'h643, 12'h643, 12'h643, 12'h642, 12'h643, 12'h643, 12'h642, 12'h643, 12'h533, 12'h532, 12'h532, 12'h532, 12'h533, 12'h532, 12'h432, 12'h433, 12'h422, 12'h422, 12'h432, 12'h433, 12'h332, 12'h322, 12'h322, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h111, 12'h111, 12'h111, 12'h333, 12'h777, 12'h777, 12'h888, 12'h999, 12'h998, 12'h999, 12'h999, 12'h988, 12'h888, 12'h888, 12'h888, 12'h887, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h877, 12'h777, 12'h777, 12'h777,
		12'h777, 12'h777, 12'h767, 12'h777, 12'h777, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h888, 12'h888, 12'h788, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h787, 12'h777, 12'h555, 12'h555, 12'h555, 12'h666, 12'h655, 12'h767, 12'h989, 12'h988, 12'h777, 12'h777, 12'h655, 12'h766, 12'h766, 12'h544, 12'h656, 12'h755, 12'h644, 12'h866, 12'h755, 12'h755, 12'h755, 12'h966, 12'h976, 12'hB76, 12'hC87, 12'hC87, 12'hC98, 12'hC98, 12'hD98, 12'hD99, 12'hEA9, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC76, 12'hC86, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'h964, 12'h955, 12'h954, 12'h964, 12'h965, 12'h954, 12'h854, 12'h854, 12'h744, 12'h743, 12'h743, 12'h643, 12'h633, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h532, 12'h432, 12'h432, 12'h532, 12'h532, 12'h422, 12'h433, 12'h432, 12'h422, 12'h422, 12'h432, 12'h333, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h111, 12'h222, 12'h121, 12'h222, 12'h211, 12'h111, 12'h222, 12'h555, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h898, 12'h989, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h787, 12'h888, 12'h878, 12'h777, 12'h777, 12'h777,
		12'h777, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h889, 12'h777, 12'h767, 12'h656, 12'h555, 12'h555, 12'h666, 12'h767, 12'h877, 12'h777, 12'h888, 12'h888, 12'h766, 12'h656, 12'h766, 12'h655, 12'h655, 12'h866, 12'h766, 12'h755, 12'h865, 12'h966, 12'h966, 12'h966, 12'hA76, 12'hB87, 12'hC98, 12'hC87, 12'hC87, 12'hC87, 12'hC98, 12'hD98, 12'hD99, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD88, 12'hD98, 12'hC87, 12'hD98, 12'hD87, 12'hD87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hD87, 12'hD87, 12'hC87, 12'hC87, 12'hD87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hB87, 12'hC87, 12'hC76, 12'hC87, 12'hB76, 12'hC86, 12'hC87, 12'hB76, 12'hB76, 12'hA65, 12'h965, 12'h965, 12'h955, 12'h954, 12'h965, 12'h964, 12'h854, 12'h854, 12'h744, 12'h743, 12'h743, 12'h643, 12'h643, 12'h633, 12'h633, 12'h633, 12'h633, 12'h532, 12'h533, 12'h533, 12'h432, 12'h533, 12'h533, 12'h422, 12'h432, 12'h432, 12'h432, 12'h432, 12'h432, 12'h322, 12'h332, 12'h332, 12'h322, 12'h222, 12'h232, 12'h222, 12'h222, 12'h232, 12'h222, 12'h211, 12'h121, 12'h222, 12'h111, 12'h111, 12'h111, 12'h444, 12'h777, 12'h888, 12'h998, 12'h999, 12'h888, 12'h988, 12'h898, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h787, 12'h877, 12'h877, 12'h787, 12'h877, 12'h777, 12'h777,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h889, 12'h888, 12'h666, 12'h666, 12'h666, 12'h656, 12'h445, 12'h545, 12'h766, 12'h777, 12'h777, 12'h877, 12'h756, 12'h655, 12'h877, 12'h977, 12'h977, 12'h966, 12'h866, 12'h976, 12'hA77, 12'hB76, 12'hB86, 12'hB87, 12'hB87, 12'hC87, 12'hB87, 12'hC87, 12'hC98, 12'hC88, 12'hC88, 12'hD98, 12'hD98, 12'hEA9, 12'hDA9, 12'hEA9, 12'hE98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD87, 12'hD98, 12'hD87, 12'hD87, 12'hD87, 12'hD87, 12'hD98, 12'hD87, 12'hD87, 12'hD87, 12'hC87, 12'hD87, 12'hD97, 12'hC87, 12'hD87, 12'hC87, 12'hC76, 12'hC87, 12'hC87, 12'hC76, 12'hC86, 12'hB76, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'h965, 12'h954, 12'h965, 12'h955, 12'h965, 12'h854, 12'h854, 12'h754, 12'h743, 12'h743, 12'h743, 12'h743, 12'h643, 12'h643, 12'h532, 12'h543, 12'h533, 12'h532, 12'h532, 12'h533, 12'h533, 12'h532, 12'h432, 12'h422, 12'h433, 12'h422, 12'h332, 12'h423, 12'h322, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h332, 12'h222, 12'h222, 12'h222, 12'h212, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h776, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h999, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h878, 12'h877, 12'h877, 12'h877, 12'h777, 12'h877,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h899, 12'h899, 12'h889, 12'h888, 12'h565, 12'h777, 12'h655, 12'h555, 12'h666, 12'h777, 12'h666, 12'h877, 12'h656, 12'h656, 12'h655, 12'h655, 12'h766, 12'h866, 12'hA88, 12'hA76, 12'h965, 12'h966, 12'hA76, 12'hC87, 12'hC87, 12'hD97, 12'hC98, 12'hC87, 12'hC87, 12'hC88, 12'hC87, 12'hD98, 12'hD98, 12'hC98, 12'hD98, 12'hD98, 12'hEA9, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD97, 12'hD87, 12'hD87, 12'hD97, 12'hC87, 12'hD98, 12'hD97, 12'hD87, 12'hD87, 12'hD87, 12'hD97, 12'hD87, 12'hD87, 12'hD87, 12'hD87, 12'hC87, 12'hD87, 12'hD87, 12'hC87, 12'hC86, 12'hC87, 12'hC87, 12'hC86, 12'hC87, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hB76, 12'hA75, 12'hA65, 12'hA65, 12'h965, 12'h965, 12'h965, 12'h955, 12'h965, 12'h954, 12'h854, 12'h854, 12'h744, 12'h744, 12'h743, 12'h743, 12'h643, 12'h643, 12'h633, 12'h532, 12'h532, 12'h533, 12'h533, 12'h532, 12'h532, 12'h422, 12'h433, 12'h432, 12'h422, 12'h322, 12'h332, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h555, 12'h877, 12'h777, 12'h888, 12'h888, 12'h998, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h787, 12'h878, 12'h877, 12'h777, 12'h878, 12'h777, 12'h877,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h787, 12'h788, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h899, 12'h899, 12'h899, 12'h899, 12'h999, 12'h877, 12'h555, 12'h556, 12'h656, 12'h666, 12'h766, 12'h667, 12'h666, 12'h766, 12'h766, 12'h666, 12'h766, 12'h655, 12'h755, 12'h976, 12'hA77, 12'hB77, 12'hA76, 12'hB77, 12'hB76, 12'hD98, 12'hD87, 12'hC87, 12'hC87, 12'hD88, 12'hC87, 12'hC98, 12'hC87, 12'hD98, 12'hD98, 12'hDA9, 12'hD98, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD97, 12'hD98, 12'hD87, 12'hD97, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD97, 12'hD87, 12'hD97, 12'hC87, 12'hC87, 12'hD87, 12'hD87, 12'hC87, 12'hC86, 12'hC87, 12'hC76, 12'hC87, 12'hC87, 12'hB87, 12'hC86, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hA75, 12'hA65, 12'h965, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'h954, 12'h955, 12'h854, 12'h854, 12'h744, 12'h743, 12'h743, 12'h643, 12'h643, 12'h633, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h532, 12'h432, 12'h433, 12'h422, 12'h432, 12'h322, 12'h332, 12'h332, 12'h322, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h333, 12'h332, 12'h222, 12'h222, 12'h121, 12'h221, 12'h222, 12'h222, 12'h111, 12'h333, 12'h777, 12'h888, 12'h999, 12'h888, 12'h999, 12'h999, 12'h988, 12'h999, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h877, 12'h878, 12'h887, 12'h877, 12'h877, 12'h777, 12'h877,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h899, 12'h899, 12'h888, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h777, 12'h555, 12'h555, 12'h455, 12'h555, 12'h888, 12'h767, 12'h656, 12'h767, 12'h767, 12'h666, 12'h877, 12'h866, 12'h866, 12'h865, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hD97, 12'hD98, 12'hD87, 12'hD87, 12'hD98, 12'hC87, 12'hD98, 12'hD98, 12'hEA9, 12'hD98, 12'hD98, 12'hEA9, 12'hEA9, 12'hE99, 12'hD99, 12'hEA9, 12'hEA9, 12'hD98, 12'hD98, 12'hE98, 12'hD98, 12'hD98, 12'hD97, 12'hE98, 12'hD98, 12'hE98, 12'hEA8, 12'hD98, 12'hD98, 12'hEA8, 12'hE98, 12'hD98, 12'hD97, 12'hC87, 12'hC87, 12'hD87, 12'hD97, 12'hC87, 12'hC97, 12'hC87, 12'hD87, 12'hC86, 12'hC86, 12'hC77, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hA65, 12'h965, 12'hA76, 12'hA65, 12'hA76, 12'hA65, 12'h965, 12'h965, 12'h954, 12'h854, 12'h854, 12'h754, 12'h743, 12'h643, 12'h643, 12'h533, 12'h643, 12'h532, 12'h532, 12'h532, 12'h533, 12'h432, 12'h433, 12'h432, 12'h422, 12'h332, 12'h422, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h666, 12'h888, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h988, 12'h988, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h877, 12'h877, 12'h878, 12'h787, 12'h877, 12'h877, 12'h877,
		12'h777, 12'h778, 12'h777, 12'h778, 12'h778, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h899, 12'h899, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h777, 12'h556, 12'h555, 12'h656, 12'h777, 12'h878, 12'h888, 12'h777, 12'h989, 12'h877, 12'h988, 12'h867, 12'h866, 12'h865, 12'h866, 12'hB87, 12'hC87, 12'hC98, 12'hD98, 12'hD98, 12'hEA9, 12'hEA9, 12'hD98, 12'hD98, 12'hDA8, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hDA9, 12'hDA9, 12'hEA9, 12'hEA9, 12'hDA9, 12'hEA9, 12'hEA9, 12'hDA9, 12'hEA9, 12'hD98, 12'hD98, 12'hD98, 12'hDA8, 12'hD97, 12'hD97, 12'hD97, 12'hD97, 12'hD98, 12'hD97, 12'hD97, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hD97, 12'hC87, 12'hD97, 12'hD98, 12'hC87, 12'hC87, 12'hC87, 12'hB76, 12'hC87, 12'hB76, 12'hB87, 12'hC87, 12'hD87, 12'hC86, 12'hB76, 12'hB76, 12'hB75, 12'hA76, 12'hA76, 12'hA76, 12'hA65, 12'hA65, 12'hA65, 12'h965, 12'h954, 12'h854, 12'h744, 12'h744, 12'h744, 12'h744, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h532, 12'h533, 12'h432, 12'h422, 12'h432, 12'h432, 12'h322, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h322, 12'h222, 12'h232, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h666, 12'h999, 12'h999, 12'h999, 12'h998, 12'h989, 12'h898, 12'h988, 12'h988, 12'h988, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h877, 12'h887, 12'h878, 12'h878, 12'h877, 12'h877, 12'h878,
		12'h878, 12'h777, 12'h878, 12'h887, 12'h788, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h999, 12'h888, 12'h667, 12'h444, 12'h555, 12'h778, 12'h777, 12'h767, 12'h888, 12'h999, 12'h888, 12'h998, 12'h766, 12'h977, 12'h866, 12'h865, 12'h965, 12'hB77, 12'hC87, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hEA9, 12'hEA9, 12'hEA9, 12'hD98, 12'hE99, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEAA, 12'hEA9, 12'hEA9, 12'hEA9, 12'hDA9, 12'hDA9, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hC98, 12'hC98, 12'hC98, 12'hC87, 12'hB87, 12'hC97, 12'hC87, 12'hC97, 12'hD98, 12'hD98, 12'hD98, 12'hC87, 12'hC87, 12'hD98, 12'hD87, 12'hC87, 12'hC87, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC76, 12'hB76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'hA76, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'h965, 12'h854, 12'h854, 12'h854, 12'h854, 12'h754, 12'h743, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h533, 12'h433, 12'h432, 12'h422, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h322, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h221, 12'h222, 12'h221, 12'h222, 12'h111, 12'h222, 12'h122, 12'h222, 12'h666, 12'h888, 12'h999, 12'h989, 12'h988, 12'h999, 12'h999, 12'h988, 12'h989, 12'h888, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h878, 12'h888, 12'h887, 12'h878, 12'h888, 12'h877, 12'h877,
		12'h888, 12'h888, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9AA, 12'h9AA, 12'h9AA, 12'h9AA, 12'h999, 12'h999, 12'h888, 12'h555, 12'h545, 12'h666, 12'h777, 12'h888, 12'h877, 12'h878, 12'h766, 12'h656, 12'h878, 12'h876, 12'h866, 12'h865, 12'hA76, 12'hC87, 12'hC87, 12'hD98, 12'hD98, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEAA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hEAA, 12'hEB9, 12'hEBA, 12'hD99, 12'hC98, 12'hC98, 12'hC98, 12'hB98, 12'hB87, 12'hA87, 12'h977, 12'h976, 12'h976, 12'h966, 12'h866, 12'h766, 12'h855, 12'h866, 12'h865, 12'hA76, 12'hA76, 12'hB87, 12'hB77, 12'hA65, 12'hC87, 12'hB86, 12'hB76, 12'hC86, 12'hC86, 12'hC86, 12'hB76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'hA65, 12'hB76, 12'hA76, 12'hA65, 12'h965, 12'h965, 12'h854, 12'h854, 12'h965, 12'h864, 12'h854, 12'h754, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h433, 12'h432, 12'h432, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h222, 12'h322, 12'h332, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h333, 12'h555, 12'h988, 12'h988, 12'h988, 12'h999, 12'h998, 12'h989, 12'h888, 12'h998, 12'h988, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h877, 12'h887, 12'h887, 12'h878, 12'h887, 12'h887,
		12'h888, 12'h888, 12'h788, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h9A9, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'h999, 12'h888, 12'h666, 12'h555, 12'h666, 12'h777, 12'h767, 12'h766, 12'h666, 12'h777, 12'h767, 12'h777, 12'h978, 12'h877, 12'h866, 12'h966, 12'hA66, 12'hB77, 12'hC87, 12'hDA8, 12'hDA9, 12'hD98, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hFA9, 12'hFBA, 12'hEBA, 12'hEB9, 12'hEBA, 12'hFBB, 12'hEBA, 12'hFBA, 12'hEB9, 12'hDA9, 12'hD98, 12'hC98, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'h976, 12'h866, 12'h755, 12'h755, 12'h855, 12'h866, 12'h755, 12'h755, 12'h755, 12'h654, 12'h644, 12'h966, 12'h855, 12'h965, 12'h855, 12'h965, 12'hA76, 12'hB76, 12'hB76, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hB86, 12'hB76, 12'hB76, 12'hA65, 12'hA65, 12'h965, 12'hA76, 12'hA75, 12'h965, 12'h965, 12'h965, 12'h965, 12'h855, 12'h854, 12'h754, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h432, 12'h533, 12'h533, 12'h543, 12'h543, 12'h532, 12'h532, 12'h433, 12'h432, 12'h332, 12'h322, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h322, 12'h332, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h555, 12'h988, 12'h888, 12'h999, 12'h999, 12'h999, 12'h988, 12'h999, 12'h999, 12'h989, 12'h888, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h878, 12'h877, 12'h888, 12'h877, 12'h887, 12'h887,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h989, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h9AA, 12'hAAA, 12'h9AA, 12'hAAA, 12'hAAA, 12'hA9A, 12'h9AA, 12'hAAA, 12'h999, 12'h777, 12'h656, 12'h666, 12'h767, 12'h888, 12'h878, 12'h878, 12'h888, 12'h988, 12'h888, 12'h877, 12'h866, 12'h865, 12'h965, 12'hA76, 12'hC87, 12'hD87, 12'hD98, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEB9, 12'hEA9, 12'hEAA, 12'hFB9, 12'hFBA, 12'hFBA, 12'hEBA, 12'hFBA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hD99, 12'hC88, 12'hB87, 12'h976, 12'hA77, 12'h977, 12'h977, 12'h976, 12'h866, 12'h976, 12'h966, 12'h966, 12'h754, 12'h654, 12'h543, 12'h755, 12'h865, 12'h644, 12'h644, 12'h543, 12'h644, 12'h754, 12'h754, 12'h754, 12'h755, 12'h854, 12'hA66, 12'hB76, 12'hC86, 12'hB76, 12'hB76, 12'hB86, 12'hC86, 12'hC87, 12'hC76, 12'hB76, 12'hB76, 12'hB76, 12'hA76, 12'hA65, 12'h965, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h755, 12'h644, 12'h533, 12'h433, 12'h433, 12'h322, 12'h221, 12'h322, 12'h222, 12'h211, 12'h321, 12'h432, 12'h432, 12'h433, 12'h432, 12'h432, 12'h432, 12'h422, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h332, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h444, 12'h777, 12'h888, 12'h999, 12'h999, 12'h988, 12'h999, 12'h998, 12'h988, 12'h999, 12'h899, 12'h988, 12'h988, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h878, 12'h887, 12'h888, 12'h878,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h999, 12'h777, 12'h666, 12'h444, 12'h666, 12'h666, 12'h777, 12'h888, 12'h988, 12'h877, 12'h877, 12'h878, 12'h866, 12'h755, 12'h865, 12'hA77, 12'hC87, 12'hD98, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEBA, 12'hEA9, 12'hFB9, 12'hEA9, 12'hEBA, 12'hFBA, 12'hEBA, 12'hEBA, 12'hEA9, 12'hFB9, 12'hDA9, 12'hD98, 12'hB87, 12'hA77, 12'hA77, 12'h976, 12'h966, 12'h966, 12'hA87, 12'hA76, 12'h965, 12'h966, 12'hA75, 12'h976, 12'h965, 12'h975, 12'h754, 12'h643, 12'h754, 12'h643, 12'h543, 12'h744, 12'h754, 12'h654, 12'h643, 12'h644, 12'h644, 12'h854, 12'h965, 12'hA76, 12'hB76, 12'hA65, 12'hA66, 12'hB76, 12'hB76, 12'hC86, 12'hB76, 12'hB75, 12'hA65, 12'hA76, 12'hA65, 12'h965, 12'h965, 12'h865, 12'h854, 12'h754, 12'h643, 12'h643, 12'h543, 12'h543, 12'h433, 12'h333, 12'h322, 12'h322, 12'h211, 12'h221, 12'h222, 12'h211, 12'h211, 12'h221, 12'h322, 12'h432, 12'h432, 12'h422, 12'h322, 12'h322, 12'h432, 12'h432, 12'h322, 12'h322, 12'h332, 12'h322, 12'h332, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h333, 12'h888, 12'h988, 12'h988, 12'h999, 12'h999, 12'h988, 12'h989, 12'h998, 12'h988, 12'h988, 12'h988, 12'h988, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h887, 12'h878, 12'h888, 12'h888,
		12'h888, 12'h888, 12'h989, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h9AA, 12'hAA9, 12'hAAA, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h888, 12'h555, 12'h545, 12'h445, 12'h666, 12'h666, 12'h888, 12'h877, 12'h877, 12'h656, 12'h766, 12'h755, 12'h755, 12'h866, 12'hA76, 12'hC87, 12'hD98, 12'hD98, 12'hEA9, 12'hEA9, 12'hEAA, 12'hEAA, 12'hEA9, 12'hEA9, 12'hFBA, 12'hFAA, 12'hEB9, 12'hFB9, 12'hEA9, 12'hEA9, 12'hD98, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hC98, 12'hB87, 12'hB87, 12'hB86, 12'hB76, 12'hB86, 12'hB76, 12'hA65, 12'hA66, 12'hA65, 12'h965, 12'h965, 12'h854, 12'h855, 12'h744, 12'h754, 12'h754, 12'h754, 12'h754, 12'h754, 12'h644, 12'h754, 12'h743, 12'h854, 12'h865, 12'h965, 12'hA65, 12'hA66, 12'hA76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA75, 12'hA65, 12'h965, 12'h965, 12'h965, 12'h854, 12'h854, 12'h754, 12'h543, 12'h533, 12'h533, 12'h433, 12'h432, 12'h332, 12'h221, 12'h221, 12'h221, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h332, 12'h332, 12'h422, 12'h433, 12'h333, 12'h322, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h777, 12'h988, 12'h988, 12'h999, 12'h999, 12'h989, 12'h999, 12'h999, 12'h989, 12'h989, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h887, 12'h888,
		12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h99A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hABA, 12'hAAA, 12'hAAA, 12'h9A9, 12'h888, 12'h555, 12'h555, 12'h544, 12'h666, 12'h778, 12'hA9A, 12'h767, 12'h766, 12'h656, 12'h655, 12'h755, 12'h765, 12'h966, 12'hB77, 12'hC87, 12'hD98, 12'hEA9, 12'hEA9, 12'hDA9, 12'hEB9, 12'hEA9, 12'hEBA, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hE98, 12'hD98, 12'hB87, 12'hB77, 12'hA77, 12'hB77, 12'hA76, 12'hB87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC87, 12'hB76, 12'hB77, 12'hB76, 12'hA76, 12'hA65, 12'h965, 12'h966, 12'h965, 12'h855, 12'h855, 12'h854, 12'h854, 12'h854, 12'h965, 12'h965, 12'h965, 12'h965, 12'h865, 12'h854, 12'h965, 12'hA76, 12'h965, 12'hA66, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA66, 12'h965, 12'h954, 12'h854, 12'h744, 12'h754, 12'h743, 12'h743, 12'h533, 12'h432, 12'h432, 12'h322, 12'h322, 12'h321, 12'h321, 12'h322, 12'h321, 12'h322, 12'h322, 12'h322, 12'h322, 12'h432, 12'h432, 12'h433, 12'h533, 12'h433, 12'h332, 12'h332, 12'h221, 12'h221, 12'h221, 12'h322, 12'h322, 12'h333, 12'h322, 12'h433, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h222, 12'h122, 12'h211, 12'h121, 12'h333, 12'h666, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h988, 12'h999, 12'h999, 12'h998, 12'h989, 12'h988, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h878, 12'h888, 12'h888, 12'h888,
		12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hABA, 12'hABA, 12'hABB, 12'hABA, 12'hABA, 12'hAAA, 12'h999, 12'h777, 12'h555, 12'h444, 12'h444, 12'h777, 12'h878, 12'h767, 12'h767, 12'h444, 12'h666, 12'h766, 12'h755, 12'h966, 12'h976, 12'hB87, 12'hC87, 12'hC98, 12'hE99, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEAA, 12'hEA9, 12'hEA9, 12'hEA8, 12'hE98, 12'hC87, 12'hC87, 12'hC87, 12'hC97, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hB87, 12'hB76, 12'hA76, 12'hA76, 12'hA66, 12'h965, 12'h965, 12'h965, 12'h854, 12'h855, 12'h854, 12'h854, 12'h854, 12'h954, 12'h955, 12'h965, 12'h965, 12'h965, 12'hA76, 12'hA65, 12'hA76, 12'hB76, 12'hC87, 12'hC86, 12'hB76, 12'hB76, 12'hA76, 12'h965, 12'h854, 12'h744, 12'h643, 12'h643, 12'h533, 12'h532, 12'h432, 12'h422, 12'h321, 12'h332, 12'h422, 12'h321, 12'h322, 12'h322, 12'h321, 12'h322, 12'h422, 12'h422, 12'h432, 12'h532, 12'h533, 12'h643, 12'h643, 12'h543, 12'h433, 12'h432, 12'h433, 12'h322, 12'h221, 12'h221, 12'h322, 12'h322, 12'h332, 12'h433, 12'h332, 12'h332, 12'h333, 12'h322, 12'h322, 12'h222, 12'h221, 12'h121, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h222, 12'h555, 12'h888, 12'h999, 12'h989, 12'h999, 12'h999, 12'h999, 12'h989, 12'h999, 12'h998, 12'h989, 12'h988, 12'h988, 12'h988, 12'h888, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888,
		12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h99A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'h999, 12'h999, 12'h656, 12'h445, 12'h545, 12'h556, 12'h656, 12'h655, 12'h655, 12'h666, 12'h877, 12'h655, 12'h755, 12'h765, 12'h865, 12'hA76, 12'hC87, 12'hC87, 12'hD98, 12'hD99, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hD98, 12'hDA9, 12'hB87, 12'hA87, 12'h966, 12'h865, 12'h865, 12'h865, 12'h865, 12'h866, 12'h755, 12'h765, 12'h765, 12'h765, 12'h765, 12'h865, 12'h865, 12'h865, 12'h755, 12'h754, 12'h644, 12'h643, 12'h643, 12'h643, 12'h643, 12'h744, 12'h754, 12'h854, 12'h854, 12'h855, 12'h854, 12'h854, 12'h854, 12'h855, 12'h965, 12'h965, 12'hA66, 12'hA76, 12'hB76, 12'hC86, 12'hC87, 12'hC87, 12'hC87, 12'hB76, 12'hA66, 12'h964, 12'h854, 12'h744, 12'h643, 12'h643, 12'h532, 12'h432, 12'h322, 12'h322, 12'h421, 12'h321, 12'h321, 12'h321, 12'h322, 12'h322, 12'h432, 12'h532, 12'h533, 12'h643, 12'h643, 12'h644, 12'h744, 12'h744, 12'h643, 12'h643, 12'h543, 12'h533, 12'h433, 12'h432, 12'h322, 12'h211, 12'h321, 12'h322, 12'h322, 12'h332, 12'h323, 12'h332, 12'h433, 12'h332, 12'h322, 12'h222, 12'h111, 12'h222, 12'h211, 12'h221, 12'h222, 12'h111, 12'h222, 12'h333, 12'h777, 12'h988, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'h989, 12'h999, 12'h989, 12'h989, 12'h988, 12'h988, 12'h988, 12'h988, 12'h888, 12'h988, 12'h888, 12'h888,
		12'h999, 12'h99A, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABA, 12'hAAA, 12'h888, 12'h666, 12'h555, 12'h555, 12'h766, 12'h666, 12'h766, 12'h767, 12'h666, 12'h655, 12'h555, 12'h756, 12'h755, 12'h966, 12'h966, 12'hC87, 12'hC87, 12'hD87, 12'hD98, 12'hEA9, 12'hD98, 12'hDA9, 12'hB87, 12'h755, 12'h332, 12'h889, 12'h545, 12'h445, 12'h222, 12'h222, 12'h333, 12'h544, 12'h755, 12'h866, 12'h976, 12'h966, 12'h976, 12'hA76, 12'h966, 12'h966, 12'h855, 12'h655, 12'h666, 12'h655, 12'h655, 12'h654, 12'h544, 12'h433, 12'h422, 12'h322, 12'h222, 12'h222, 12'h222, 12'h322, 12'h422, 12'h533, 12'h643, 12'h744, 12'h854, 12'h955, 12'hA65, 12'hA76, 12'hB76, 12'hB76, 12'hC76, 12'hC76, 12'hC87, 12'hB76, 12'hA66, 12'h854, 12'h754, 12'h643, 12'h533, 12'h432, 12'h321, 12'h321, 12'h322, 12'h321, 12'h321, 12'h322, 12'h432, 12'h433, 12'h533, 12'h643, 12'h644, 12'h754, 12'h754, 12'h754, 12'h754, 12'h854, 12'h754, 12'h754, 12'h743, 12'h643, 12'h643, 12'h643, 12'h533, 12'h432, 12'h432, 12'h322, 12'h221, 12'h222, 12'h322, 12'h322, 12'h332, 12'h433, 12'h332, 12'h323, 12'h332, 12'h222, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h333, 12'h777, 12'h988, 12'h999, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'hA99, 12'h999, 12'h998, 12'h988, 12'h988, 12'h989, 12'h988, 12'h989, 12'h988, 12'h988, 12'h989, 12'h888, 12'h888,
		12'h999, 12'h99A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hABB, 12'hBBA, 12'hABB, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABA, 12'h888, 12'h766, 12'h444, 12'h656, 12'h666, 12'h555, 12'h666, 12'h767, 12'h666, 12'h877, 12'h655, 12'h655, 12'h755, 12'h866, 12'h965, 12'hA76, 12'hB76, 12'hB87, 12'hC87, 12'hD98, 12'hA76, 12'h544, 12'h222, 12'h777, 12'h333, 12'hA9A, 12'h445, 12'h445, 12'h223, 12'h333, 12'h645, 12'hA76, 12'hA76, 12'hB76, 12'hA76, 12'hA76, 12'h976, 12'h966, 12'h644, 12'h644, 12'h755, 12'h866, 12'h866, 12'h866, 12'h866, 12'h866, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h432, 12'h644, 12'h644, 12'h533, 12'h433, 12'h432, 12'h322, 12'h422, 12'h533, 12'h955, 12'hA65, 12'hB76, 12'hB76, 12'hB77, 12'hC87, 12'hB76, 12'hA76, 12'h966, 12'h854, 12'h643, 12'h533, 12'h322, 12'h322, 12'h321, 12'h221, 12'h221, 12'h321, 12'h432, 12'h433, 12'h543, 12'h643, 12'h744, 12'h744, 12'h654, 12'h744, 12'h744, 12'h754, 12'h754, 12'h854, 12'h854, 12'h754, 12'h744, 12'h754, 12'h643, 12'h533, 12'h432, 12'h432, 12'h322, 12'h322, 12'h321, 12'h221, 12'h222, 12'h322, 12'h322, 12'h332, 12'h322, 12'h333, 12'h332, 12'h222, 12'h211, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h444, 12'h877, 12'h888, 12'hA99, 12'hAAA, 12'hA9A, 12'h9A9, 12'hA9A, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h989, 12'h998, 12'h999, 12'h999, 12'h999, 12'h988, 12'h999, 12'h999, 12'h988, 12'h988,
		12'h999, 12'h999, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hABA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABA, 12'h889, 12'h666, 12'h545, 12'h444, 12'h656, 12'h555, 12'h444, 12'h555, 12'h767, 12'h544, 12'h545, 12'h544, 12'h644, 12'h644, 12'h755, 12'h854, 12'h955, 12'h754, 12'h644, 12'h434, 12'h334, 12'h433, 12'h223, 12'h444, 12'h222, 12'hAAB, 12'h334, 12'h444, 12'h333, 12'h333, 12'h976, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h976, 12'h866, 12'h655, 12'h655, 12'h866, 12'h966, 12'hA77, 12'hB88, 12'hA77, 12'h865, 12'h755, 12'h754, 12'h533, 12'h433, 12'h543, 12'h533, 12'h533, 12'h422, 12'h533, 12'h644, 12'h744, 12'h744, 12'h754, 12'h755, 12'h754, 12'h443, 12'h422, 12'h955, 12'hB76, 12'hB76, 12'hB77, 12'hC87, 12'hB86, 12'hA65, 12'h854, 12'h643, 12'h432, 12'h322, 12'h221, 12'h211, 12'h211, 12'h322, 12'h432, 12'h322, 12'h321, 12'h211, 12'h221, 12'h221, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h221, 12'h222, 12'h221, 12'h222, 12'h221, 12'h321, 12'h222, 12'h221, 12'h322, 12'h322, 12'h221, 12'h221, 12'h222, 12'h322, 12'h322, 12'h332, 12'h322, 12'h433, 12'h332, 12'h222, 12'h221, 12'h121, 12'h111, 12'h111, 12'h222, 12'h222, 12'h111, 12'h444, 12'h666, 12'h888, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'h999, 12'h999, 12'hA99, 12'hA89, 12'h989, 12'h999, 12'h988, 12'h988, 12'h999, 12'h999, 12'h988, 12'h999, 12'h998, 12'h999,
		12'h999, 12'hAAA, 12'hAAA, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABA, 12'hBBB, 12'hBAA, 12'h877, 12'h666, 12'h444, 12'h555, 12'h544, 12'h545, 12'h434, 12'h444, 12'h555, 12'h556, 12'h555, 12'h555, 12'h333, 12'h333, 12'h433, 12'h433, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h533, 12'h533, 12'h643, 12'h755, 12'h644, 12'h433, 12'h322, 12'h544, 12'hA76, 12'hB77, 12'hA77, 12'hA77, 12'h976, 12'h876, 12'h766, 12'h866, 12'h866, 12'h965, 12'h855, 12'h645, 12'h433, 12'h545, 12'h545, 12'h444, 12'h323, 12'h322, 12'h333, 12'h433, 12'h433, 12'h433, 12'h432, 12'h422, 12'h433, 12'h644, 12'h643, 12'h744, 12'h855, 12'h966, 12'hA76, 12'hA77, 12'h333, 12'h433, 12'h643, 12'h643, 12'h643, 12'h543, 12'h533, 12'h433, 12'h432, 12'h322, 12'h321, 12'h221, 12'h432, 12'h322, 12'h432, 12'h322, 12'h323, 12'h322, 12'h433, 12'h433, 12'h543, 12'h755, 12'h965, 12'h865, 12'h855, 12'h754, 12'h744, 12'h644, 12'h533, 12'h432, 12'h432, 12'h533, 12'h433, 12'h433, 12'h432, 12'h322, 12'h322, 12'h222, 12'h222, 12'h322, 12'h222, 12'h221, 12'h221, 12'h222, 12'h322, 12'h322, 12'h322, 12'h222, 12'h211, 12'h111, 12'h222, 12'h222, 12'h222, 12'h221, 12'h111, 12'h222, 12'h666, 12'h999, 12'hA99, 12'hAAA, 12'hA99, 12'hA9A, 12'hA9A, 12'hA99, 12'hA99, 12'h999, 12'h999, 12'hA99, 12'h989, 12'h999, 12'h989, 12'h999, 12'h988, 12'h999, 12'h988, 12'h999, 12'h999,
		12'h99A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hABB, 12'hBBB, 12'hBBB, 12'hAAA, 12'h887, 12'h666, 12'h655, 12'h545, 12'h444, 12'h444, 12'h555, 12'h545, 12'h544, 12'h555, 12'h777, 12'h877, 12'h544, 12'h222, 12'h222, 12'h322, 12'h555, 12'h767, 12'hA87, 12'hB88, 12'hB76, 12'hA76, 12'hB76, 12'hA76, 12'hA66, 12'hA75, 12'hA65, 12'h855, 12'h333, 12'h755, 12'hA66, 12'hB87, 12'hB87, 12'hA87, 12'h987, 12'h987, 12'h977, 12'h976, 12'h754, 12'h544, 12'h656, 12'h767, 12'h445, 12'hCCC, 12'h556, 12'h344, 12'h433, 12'h434, 12'h656, 12'h877, 12'h533, 12'h322, 12'h433, 12'h433, 12'h432, 12'h433, 12'h533, 12'h644, 12'h855, 12'h976, 12'hA77, 12'hB88, 12'h877, 12'h111, 12'h221, 12'h311, 12'h433, 12'h543, 12'h533, 12'h322, 12'h211, 12'h111, 12'h111, 12'h555, 12'h111, 12'h555, 12'h322, 12'h333, 12'h333, 12'h322, 12'h333, 12'h655, 12'h866, 12'h966, 12'h977, 12'h966, 12'h966, 12'h854, 12'h643, 12'h643, 12'h533, 12'h433, 12'h432, 12'h322, 12'h322, 12'h432, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h333, 12'h544, 12'h545, 12'h555, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h221, 12'h111, 12'h121, 12'h112, 12'h111, 12'h222, 12'h222, 12'h777, 12'h999, 12'hA9A, 12'hAAA, 12'hAA9, 12'hA9A, 12'hA9A, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h989, 12'h999, 12'h989, 12'h988, 12'h999, 12'h999,
		12'h9AA, 12'hA99, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBA, 12'hCCB, 12'hECC, 12'hEBB, 12'hDA9, 12'hB87, 12'h855, 12'h644, 12'h444, 12'h555, 12'h766, 12'h666, 12'h655, 12'h444, 12'h333, 12'h655, 12'h544, 12'h656, 12'h977, 12'hCBA, 12'hECC, 12'hECB, 12'hEAA, 12'hEA9, 12'hEA9, 12'hD98, 12'hD98, 12'hD98, 12'hC87, 12'hB77, 12'hB87, 12'hB87, 12'h544, 12'h966, 12'hA77, 12'hB87, 12'hB98, 12'hB88, 12'hA88, 12'hA87, 12'h876, 12'h755, 12'h755, 12'h856, 12'hA88, 12'hBAA, 12'h545, 12'h434, 12'h433, 12'h433, 12'h433, 12'h655, 12'hA9A, 12'hCAA, 12'h967, 12'h544, 12'h433, 12'h533, 12'h433, 12'h433, 12'h533, 12'h755, 12'h967, 12'hA76, 12'hA66, 12'hB88, 12'h666, 12'h543, 12'h643, 12'h965, 12'hC87, 12'hC87, 12'hA75, 12'h854, 12'h533, 12'h321, 12'h210, 12'h322, 12'h100, 12'h655, 12'h222, 12'h333, 12'h333, 12'h433, 12'h644, 12'h755, 12'h856, 12'h645, 12'h644, 12'h544, 12'h333, 12'h333, 12'h323, 12'h332, 12'h422, 12'h432, 12'h433, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h322, 12'h332, 12'h433, 12'h222, 12'h544, 12'h777, 12'h222, 12'h111, 12'h121, 12'h111, 12'h221, 12'h111, 12'h111, 12'h222, 12'h111, 12'h121, 12'h222, 12'h333, 12'h777, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA99, 12'hAAA, 12'hA9A, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'h989, 12'hA99, 12'h989, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBAA, 12'h954, 12'hA65, 12'hC87, 12'hEAA, 12'hEA8, 12'hC87, 12'hA66, 12'h855, 12'h544, 12'h766, 12'h545, 12'h433, 12'h434, 12'h434, 12'h544, 12'h766, 12'hA88, 12'hC98, 12'hEBA, 12'hEBA, 12'hFBA, 12'hEA9, 12'hEA9, 12'hEA8, 12'hDA8, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'h543, 12'hB87, 12'hC87, 12'hC98, 12'hC98, 12'hB98, 12'hB88, 12'hA88, 12'hA87, 12'hA77, 12'hA77, 12'hB87, 12'hB88, 12'hB77, 12'hA88, 12'h766, 12'h544, 12'h433, 12'h534, 12'h656, 12'hB99, 12'hB98, 12'h966, 12'h755, 12'h744, 12'h644, 12'h533, 12'h533, 12'h534, 12'h877, 12'hA77, 12'hA77, 12'hA76, 12'hCAA, 12'h444, 12'h422, 12'h854, 12'hD87, 12'hD97, 12'hD87, 12'hB76, 12'h964, 12'h743, 12'h432, 12'h210, 12'h322, 12'h111, 12'h655, 12'h322, 12'h433, 12'h544, 12'h544, 12'h544, 12'h433, 12'h433, 12'h444, 12'h334, 12'hDCD, 12'h667, 12'h334, 12'h333, 12'h333, 12'h333, 12'h322, 12'h222, 12'h322, 12'h332, 12'h322, 12'h322, 12'h222, 12'h322, 12'h332, 12'h332, 12'h433, 12'h433, 12'h222, 12'h444, 12'h889, 12'h544, 12'h121, 12'h111, 12'h111, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h666, 12'h767, 12'hA99, 12'hAAA, 12'hBAA, 12'hA9A, 12'hAAA, 12'hAA9, 12'hAAA, 12'hA9A, 12'hA9A, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'h999, 12'hA99, 12'h999, 12'hA99, 12'hA99, 12'hA99,
		12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hABB, 12'hBBB, 12'hBBB, 12'hABB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBBB, 12'hBCC, 12'hBCB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hBBA, 12'h843, 12'h843, 12'h943, 12'hA65, 12'hC87, 12'hD99, 12'hC87, 12'h966, 12'h988, 12'h877, 12'h666, 12'h444, 12'h444, 12'h434, 12'h655, 12'hA87, 12'hD98, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA8, 12'hE98, 12'hEA8, 12'hE98, 12'h654, 12'hB88, 12'hD98, 12'hD99, 12'hDA9, 12'hCA9, 12'hC99, 12'hC99, 12'hC88, 12'hB87, 12'hC88, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hA87, 12'hB88, 12'h966, 12'h755, 12'h754, 12'h644, 12'h644, 12'h643, 12'h543, 12'h533, 12'h544, 12'h433, 12'h655, 12'h655, 12'h766, 12'h966, 12'hA76, 12'hA77, 12'hBAA, 12'h211, 12'h533, 12'hA76, 12'hFA8, 12'hFA9, 12'hE98, 12'hD86, 12'hB65, 12'h854, 12'h533, 12'h221, 12'h221, 12'h111, 12'h544, 12'h433, 12'h545, 12'h544, 12'h433, 12'h433, 12'h545, 12'h988, 12'hA99, 12'h445, 12'h544, 12'h333, 12'h333, 12'h333, 12'h444, 12'h656, 12'h555, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h322, 12'h332, 12'h322, 12'h432, 12'h433, 12'h433, 12'h323, 12'h444, 12'h889, 12'h666, 12'h211, 12'h221, 12'h221, 12'h222, 12'h121, 12'h111, 12'h111, 12'h221, 12'h222, 12'h445, 12'h777, 12'h888, 12'hAAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA9A, 12'hA9A, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'h999, 12'hA99, 12'hAAA, 12'hAAA,
		12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hA87, 12'hA54, 12'hB55, 12'hB75, 12'hC76, 12'hC86, 12'hD98, 12'hC98, 12'hB87, 12'h966, 12'h866, 12'h544, 12'h444, 12'h545, 12'h766, 12'hC98, 12'hD98, 12'hD98, 12'hEA9, 12'hEA9, 12'hDA8, 12'hEA9, 12'hEA8, 12'hE99, 12'hEA9, 12'hEA9, 12'hEA8, 12'hEA9, 12'hEA8, 12'hEA9, 12'hEA8, 12'h965, 12'hA77, 12'hEA9, 12'hDA9, 12'hEA9, 12'hDA9, 12'hDA9, 12'hDA8, 12'hD98, 12'hC87, 12'hC88, 12'hB87, 12'hB88, 12'hB88, 12'hA77, 12'hA77, 12'hA76, 12'h966, 12'h855, 12'h754, 12'h644, 12'h644, 12'h644, 12'h533, 12'h534, 12'h544, 12'h544, 12'h644, 12'h755, 12'h866, 12'h977, 12'h977, 12'hA88, 12'h888, 12'h322, 12'h744, 12'hE98, 12'hFB9, 12'hFB9, 12'hFB9, 12'hE97, 12'hC86, 12'hA65, 12'h633, 12'h322, 12'h321, 12'h110, 12'h444, 12'h333, 12'h434, 12'h333, 12'h433, 12'h544, 12'h644, 12'h755, 12'h987, 12'h767, 12'h666, 12'h544, 12'h433, 12'h433, 12'h544, 12'h654, 12'h644, 12'h433, 12'h322, 12'h222, 12'h222, 12'h222, 12'h322, 12'h422, 12'h432, 12'h433, 12'h433, 12'h433, 12'h322, 12'h434, 12'h888, 12'h665, 12'h221, 12'h322, 12'h221, 12'h111, 12'h221, 12'h221, 12'h111, 12'h221, 12'h333, 12'h444, 12'h777, 12'hAAA, 12'hAAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA9A, 12'hA9A, 12'hA99, 12'hA99, 12'hA99, 12'hA9A, 12'hAAA, 12'hAA9, 12'hAA9,
		12'hAAA, 12'hABB, 12'hBBB, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBCC, 12'hCCB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCAA, 12'hC75, 12'hC76, 12'hC76, 12'hD86, 12'hD87, 12'hC86, 12'hC88, 12'hC87, 12'hB77, 12'h866, 12'h755, 12'h644, 12'h644, 12'hA77, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEB9, 12'hEA8, 12'hEA9, 12'hEA8, 12'hEA8, 12'hC86, 12'h765, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA8, 12'hE98, 12'hD98, 12'hD87, 12'hC87, 12'hB87, 12'hB77, 12'hA76, 12'hA66, 12'h965, 12'h965, 12'h865, 12'h855, 12'h855, 12'h754, 12'h744, 12'h644, 12'h644, 12'h744, 12'h755, 12'h755, 12'h856, 12'h966, 12'h976, 12'hA77, 12'h766, 12'hBAA, 12'h443, 12'h322, 12'hA65, 12'hFA9, 12'hFCA, 12'hFB9, 12'hFB9, 12'hE97, 12'hD86, 12'hB75, 12'h843, 12'h322, 12'h222, 12'h111, 12'h333, 12'h322, 12'h544, 12'h544, 12'h544, 12'h655, 12'h655, 12'h755, 12'h765, 12'h866, 12'h755, 12'h765, 12'h754, 12'h744, 12'h643, 12'h533, 12'h643, 12'h543, 12'h533, 12'h432, 12'h322, 12'h322, 12'h322, 12'h332, 12'h432, 12'h433, 12'h533, 12'h433, 12'h444, 12'h888, 12'hAAA, 12'h777, 12'h322, 12'h333, 12'h111, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h444, 12'h667, 12'h999, 12'hBBB, 12'hBBB, 12'hBAA, 12'hBBB, 12'hBBA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA9A, 12'hA9A, 12'hAAA, 12'hA99, 12'hAA9, 12'hA99, 12'hA99,
		12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBC, 12'hBBB, 12'hCCC, 12'hBCC, 12'hCCB, 12'hBCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hC75, 12'hC75, 12'hD86, 12'hD86, 12'hE97, 12'hE98, 12'hC87, 12'hD97, 12'hD98, 12'hC87, 12'hA76, 12'h855, 12'h654, 12'hA77, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEB9, 12'hFA9, 12'hEA9, 12'hFB9, 12'hEA9, 12'hEA8, 12'hEA8, 12'h644, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA8, 12'hEA8, 12'hE98, 12'hD98, 12'hD88, 12'hC87, 12'hC87, 12'hB77, 12'hA77, 12'hA66, 12'hA66, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h966, 12'hA77, 12'hA77, 12'h866, 12'h877, 12'hA99, 12'h221, 12'h743, 12'hD97, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hF98, 12'hE86, 12'hC75, 12'h854, 12'h432, 12'h322, 12'h111, 12'h221, 12'h433, 12'h433, 12'h533, 12'h544, 12'h644, 12'h544, 12'h655, 12'h755, 12'h755, 12'h755, 12'h754, 12'h644, 12'h643, 12'h643, 12'h543, 12'h533, 12'h533, 12'h433, 12'h432, 12'h433, 12'h433, 12'h432, 12'h432, 12'h433, 12'h533, 12'h543, 12'h433, 12'h556, 12'h999, 12'hBBC, 12'h888, 12'h333, 12'h332, 12'h222, 12'h221, 12'h222, 12'h222, 12'h444, 12'h444, 12'h444, 12'h888, 12'hBAA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBAA, 12'hAAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA99, 12'hAAA, 12'hAAA, 12'hA99, 12'hA99, 12'hA99, 12'hA99,
		12'hABA, 12'hBBA, 12'hABB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCA8, 12'hD86, 12'hD86, 12'hD87, 12'hFB9, 12'hFBA, 12'hEA8, 12'hC86, 12'hD87, 12'hD87, 12'hC87, 12'hA76, 12'h976, 12'hB87, 12'hD99, 12'hD98, 12'hDA8, 12'hD98, 12'hE98, 12'hDA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hEA9, 12'h754, 12'hB87, 12'hE98, 12'hEA9, 12'hFB9, 12'hFA9, 12'hEA9, 12'hEA9, 12'hEA8, 12'hE98, 12'hE98, 12'hD98, 12'hD88, 12'hD88, 12'hC87, 12'hC87, 12'hB77, 12'hB76, 12'hA66, 12'h966, 12'h965, 12'h965, 12'h966, 12'h966, 12'h966, 12'h966, 12'hA76, 12'hA77, 12'h966, 12'h877, 12'hAAA, 12'h333, 12'h633, 12'hC87, 12'hFA9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFA8, 12'hE97, 12'hC76, 12'h954, 12'h532, 12'h221, 12'h222, 12'h110, 12'h433, 12'h433, 12'h543, 12'h644, 12'h644, 12'h744, 12'h744, 12'h754, 12'h744, 12'h644, 12'h644, 12'h643, 12'h643, 12'h533, 12'h533, 12'h543, 12'h533, 12'h533, 12'h543, 12'h643, 12'h543, 12'h433, 12'h433, 12'h433, 12'h533, 12'h543, 12'h433, 12'h545, 12'hA9A, 12'hEDE, 12'h555, 12'h432, 12'h322, 12'h322, 12'h222, 12'h121, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h433, 12'h544, 12'h887, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABB, 12'hBBA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hA9A, 12'hAAA, 12'hA99, 12'hA9A, 12'hAAA,
		12'hABA, 12'hBBB, 12'hABB, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hDBA, 12'hD98, 12'hE98, 12'hF98, 12'hFCA, 12'hFCB, 12'hFBB, 12'hE98, 12'hD86, 12'hD87, 12'hD87, 12'hB76, 12'h976, 12'hC98, 12'hD99, 12'hDA8, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEBA, 12'hEBA, 12'hFCA, 12'hFCA, 12'hFCA, 12'hFCB, 12'hFCB, 12'hFBA, 12'hEBA, 12'h544, 12'hB87, 12'hEA9, 12'hEA9, 12'hFA9, 12'hEA8, 12'hEA8, 12'hE98, 12'hE98, 12'hEA9, 12'hEA9, 12'hE98, 12'hE98, 12'hD98, 12'hD88, 12'hC87, 12'hB77, 12'hB76, 12'hB66, 12'hA66, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hC87, 12'hB87, 12'hB76, 12'hA66, 12'hBA9, 12'h433, 12'h633, 12'hB77, 12'hFA9, 12'hFBA, 12'hFB9, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFA8, 12'hE97, 12'hD76, 12'hA54, 12'h643, 12'h322, 12'h221, 12'h111, 12'h322, 12'h433, 12'h533, 12'h644, 12'h755, 12'h755, 12'h855, 12'h855, 12'h754, 12'h744, 12'h754, 12'h744, 12'h754, 12'h744, 12'h744, 12'h744, 12'h754, 12'h744, 12'h754, 12'h644, 12'h644, 12'h543, 12'h433, 12'h533, 12'h533, 12'h444, 12'h444, 12'h555, 12'hBAB, 12'hEDE, 12'h322, 12'h332, 12'h332, 12'h322, 12'h222, 12'h111, 12'h211, 12'h221, 12'h322, 12'h322, 12'h432, 12'h332, 12'h322, 12'h222, 12'hBAA, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hBAA, 12'hAAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hDDC, 12'hDDC, 12'hE98, 12'hEA9, 12'hFA9, 12'hFBA, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFCB, 12'hC76, 12'hC86, 12'hC86, 12'hB76, 12'hA77, 12'hC88, 12'hD98, 12'hD98, 12'hE98, 12'hD98, 12'hEA9, 12'hDA8, 12'hEA9, 12'hEA9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFCA, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFBA, 12'hFBA, 12'hEA9, 12'h965, 12'h754, 12'h866, 12'hC97, 12'hEA8, 12'hEA8, 12'hE98, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hE98, 12'hD98, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC76, 12'hB76, 12'hC77, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC87, 12'hB88, 12'h544, 12'h533, 12'hA65, 12'hFA8, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA9, 12'hFB9, 12'hFA9, 12'hF98, 12'hF97, 12'hD86, 12'hA65, 12'h743, 12'h532, 12'h322, 12'h221, 12'h111, 12'h533, 12'h643, 12'h643, 12'h643, 12'h754, 12'h865, 12'h965, 12'h966, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h744, 12'h754, 12'h754, 12'h754, 12'h744, 12'h644, 12'h543, 12'h533, 12'h543, 12'h543, 12'h533, 12'h444, 12'h656, 12'hDCD, 12'h888, 12'h333, 12'h332, 12'h322, 12'h322, 12'h222, 12'h221, 12'h221, 12'h322, 12'h432, 12'h432, 12'h322, 12'h221, 12'h211, 12'h222, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBAA, 12'hBAB, 12'hAAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDC, 12'hDDD, 12'hEBB, 12'hD76, 12'hE98, 12'hFA8, 12'hFCA, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFCB, 12'hE98, 12'hB75, 12'hB76, 12'hA66, 12'hA77, 12'hC98, 12'hD98, 12'hD98, 12'hEA9, 12'hD99, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEB9, 12'hEB9, 12'hFBA, 12'hFBA, 12'hFCB, 12'hEBB, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFBA, 12'hEB9, 12'hD98, 12'hD97, 12'hC76, 12'h854, 12'h744, 12'h644, 12'h755, 12'hA76, 12'hB98, 12'hD99, 12'hDA9, 12'hD98, 12'hD98, 12'hD88, 12'hC76, 12'hC87, 12'hC87, 12'hD87, 12'hC87, 12'hD97, 12'hD98, 12'hD98, 12'hD98, 12'hC88, 12'hB88, 12'h977, 12'h543, 12'h633, 12'hA66, 12'hE98, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hF97, 12'hF87, 12'hD76, 12'hA65, 12'h843, 12'h533, 12'h422, 12'h322, 12'h321, 12'h322, 12'h644, 12'h744, 12'h744, 12'h744, 12'h744, 12'h854, 12'h855, 12'h855, 12'h955, 12'h854, 12'h854, 12'h844, 12'h754, 12'h854, 12'h743, 12'h854, 12'h854, 12'h754, 12'h753, 12'h643, 12'h533, 12'h543, 12'h543, 12'h533, 12'h544, 12'h767, 12'hEEE, 12'h443, 12'h332, 12'h322, 12'h322, 12'h332, 12'h332, 12'h222, 12'h322, 12'h322, 12'h332, 12'h322, 12'h221, 12'h211, 12'h211, 12'h666, 12'hCCB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hABA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDAA, 12'hC76, 12'hD98, 12'hFA8, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hE86, 12'hA64, 12'h966, 12'hA76, 12'hC98, 12'hD98, 12'hD98, 12'hDA9, 12'hDA8, 12'hDA8, 12'hD98, 12'hEA9, 12'hFB9, 12'hEA9, 12'hEB9, 12'hEBA, 12'hFBA, 12'hFBA, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFCA, 12'hFCA, 12'hFBA, 12'hFB9, 12'hFA8, 12'hE98, 12'hE97, 12'hD86, 12'hC86, 12'hC76, 12'hB75, 12'h954, 12'h843, 12'h743, 12'h754, 12'h754, 12'h754, 12'h755, 12'h755, 12'h754, 12'h754, 12'h744, 12'h744, 12'h644, 12'h744, 12'h643, 12'h643, 12'h533, 12'h532, 12'h643, 12'hA65, 12'hD88, 12'hE98, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hFA8, 12'hF97, 12'hF97, 12'hE87, 12'hD86, 12'hB65, 12'h854, 12'h743, 12'h533, 12'h432, 12'h422, 12'h321, 12'h432, 12'h643, 12'h754, 12'h754, 12'h744, 12'h853, 12'h743, 12'h854, 12'h854, 12'h854, 12'h844, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h744, 12'h643, 12'h644, 12'h544, 12'h544, 12'h545, 12'hBBB, 12'h766, 12'h433, 12'h332, 12'h332, 12'h322, 12'h322, 12'h332, 12'h221, 12'h321, 12'h322, 12'h321, 12'h221, 12'h221, 12'h311, 12'h322, 12'hBBB, 12'hCCB, 12'hCCC, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hAAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDC, 12'hDDD, 12'hEA9, 12'hC76, 12'hD99, 12'hFA9, 12'hFA8, 12'hF97, 12'hF87, 12'hE86, 12'hD75, 12'hA54, 12'h743, 12'hB77, 12'hB87, 12'hC98, 12'hDA9, 12'hD98, 12'hDA9, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hFB9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hEBA, 12'hFBA, 12'hFCA, 12'hFBB, 12'hFBA, 12'hFCB, 12'hFBA, 12'hFB9, 12'hFA9, 12'hFA8, 12'hD98, 12'hFA8, 12'hE98, 12'hE97, 12'hE97, 12'hD87, 12'hB76, 12'hB76, 12'hB76, 12'hB65, 12'hB65, 12'hA65, 12'hB65, 12'hB65, 12'hA65, 12'hA65, 12'hB65, 12'hA65, 12'hB65, 12'hB66, 12'hB76, 12'hC87, 12'hD98, 12'hE98, 12'hE99, 12'hEA9, 12'hFA8, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hFA8, 12'hF98, 12'hFA8, 12'hF97, 12'hE97, 12'hD86, 12'hC76, 12'hA65, 12'h854, 12'h743, 12'h533, 12'h432, 12'h432, 12'h321, 12'h211, 12'h221, 12'h432, 12'h533, 12'h744, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h964, 12'h965, 12'h964, 12'h954, 12'h854, 12'h854, 12'h754, 12'h755, 12'h766, 12'h666, 12'h545, 12'h332, 12'h333, 12'h332, 12'h323, 12'h333, 12'h322, 12'h322, 12'h333, 12'h222, 12'h321, 12'h322, 12'h221, 12'h321, 12'h221, 12'h321, 12'h766, 12'hCCC, 12'hCCC, 12'hCBB, 12'hBBB, 12'hCCB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hAAA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA, 12'hAAA,
		12'hBBB, 12'hBCB, 12'hBCB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDD, 12'hDCC, 12'hE97, 12'hC76, 12'hE98, 12'hFA9, 12'hE97, 12'hD86, 12'hD76, 12'hC75, 12'hB65, 12'hA54, 12'h954, 12'hC98, 12'hB98, 12'hC98, 12'hC98, 12'hD98, 12'hD98, 12'hD98, 12'hDA8, 12'hD98, 12'hEA9, 12'hEA9, 12'hEB9, 12'hEA9, 12'hEAA, 12'hEBA, 12'hFBA, 12'hEB9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hFA8, 12'hEA8, 12'hE97, 12'hE97, 12'hD87, 12'hE97, 12'hD97, 12'hD87, 12'hE98, 12'hE98, 12'hE98, 12'hD97, 12'hD97, 12'hD97, 12'hE97, 12'hE98, 12'hD98, 12'hE98, 12'hEA9, 12'hFA9, 12'hEAA, 12'hEA9, 12'hE98, 12'hE98, 12'hF98, 12'hF98, 12'hFA8, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hF97, 12'hF97, 12'hE97, 12'hD86, 12'hD86, 12'hB65, 12'hA65, 12'h854, 12'h643, 12'h432, 12'h432, 12'h533, 12'h533, 12'h532, 12'h421, 12'h311, 12'h211, 12'h221, 12'h321, 12'h322, 12'h432, 12'h432, 12'h533, 12'h533, 12'h543, 12'h643, 12'h644, 12'h544, 12'h544, 12'h544, 12'h433, 12'h332, 12'h322, 12'h322, 12'h321, 12'h322, 12'h433, 12'h432, 12'h322, 12'h432, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h221, 12'h322, 12'h221, 12'h311, 12'h221, 12'h322, 12'hAAA, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCCB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBBA, 12'hBAA, 12'hBAA, 12'hAAA, 12'hBAA, 12'hAAA, 12'hAAA,
		12'hBCB, 12'hBBB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCB, 12'hBBB, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDCC, 12'hE98, 12'hC76, 12'hE98, 12'hFA9, 12'hE87, 12'hD76, 12'hC75, 12'hB65, 12'hA64, 12'hA54, 12'hA65, 12'hC87, 12'hB88, 12'hC99, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEB9, 12'hEA9, 12'hEA9, 12'hEBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFCA, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hE98, 12'hF98, 12'hE98, 12'hE97, 12'hE97, 12'hE98, 12'hE98, 12'hE98, 12'hE98, 12'hE97, 12'hE97, 12'hE98, 12'hE97, 12'hE98, 12'hE98, 12'hEA8, 12'hEA9, 12'hEA9, 12'hE99, 12'hD98, 12'hD87, 12'hE87, 12'hE97, 12'hE98, 12'hFA8, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFA8, 12'hFA8, 12'hF98, 12'hF97, 12'hE87, 12'hD87, 12'hC75, 12'hB65, 12'h965, 12'h854, 12'h643, 12'h432, 12'h533, 12'h533, 12'h643, 12'h743, 12'h643, 12'h643, 12'h643, 12'h632, 12'h632, 12'h532, 12'h532, 12'h532, 12'h633, 12'h633, 12'h633, 12'h643, 12'h643, 12'h743, 12'h643, 12'h643, 12'h643, 12'h643, 12'h532, 12'h432, 12'h432, 12'h432, 12'h322, 12'h322, 12'h333, 12'h332, 12'h333, 12'h322, 12'h332, 12'h222, 12'h321, 12'h322, 12'h221, 12'h321, 12'h321, 12'h433, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hBBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBAB, 12'hBBB, 12'hBAA, 12'hBAB, 12'hBAA, 12'hBAA, 12'hAAA, 12'hAAA,
		12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hBCC, 12'hBCB, 12'hCCC, 12'hCBC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDD, 12'hDCC, 12'hD98, 12'hC76, 12'hE98, 12'hFBA, 12'hE87, 12'hC75, 12'hC65, 12'hB65, 12'hB65, 12'hB75, 12'hB76, 12'hC87, 12'hC99, 12'hC98, 12'hC98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hFBA, 12'hFA9, 12'hEB9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hF98, 12'hFA8, 12'hFA8, 12'hFA8, 12'hE98, 12'hEA8, 12'hE98, 12'hE97, 12'hE97, 12'hD87, 12'hD87, 12'hD87, 12'hD87, 12'hD98, 12'hD98, 12'hD87, 12'hD87, 12'hD87, 12'hE98, 12'hFA8, 12'hFA8, 12'hFB9, 12'hFB9, 12'hFCA, 12'hFCA, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFA8, 12'hFA8, 12'hF98, 12'hE97, 12'hD86, 12'hC76, 12'hA65, 12'h954, 12'h854, 12'h643, 12'h533, 12'h432, 12'h533, 12'h753, 12'h843, 12'h854, 12'h954, 12'h854, 12'h854, 12'h854, 12'h843, 12'h754, 12'h743, 12'h743, 12'h753, 12'h743, 12'h743, 12'h743, 12'h743, 12'h643, 12'h633, 12'h533, 12'h532, 12'h432, 12'h432, 12'h332, 12'h332, 12'h433, 12'h422, 12'h333, 12'h323, 12'h332, 12'h332, 12'h222, 12'h321, 12'h322, 12'h221, 12'h321, 12'h322, 12'h877, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBAB, 12'hBBB, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBAA, 12'hAAA, 12'hABA, 12'hBAA,
		12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDAA, 12'hD88, 12'hE98, 12'hFBA, 12'hE97, 12'hD76, 12'hC65, 12'hB65, 12'hB65, 12'hC75, 12'hC76, 12'hB77, 12'hC98, 12'hC98, 12'hC98, 12'hD98, 12'hD98, 12'hC97, 12'hD98, 12'hD98, 12'hD98, 12'hEA8, 12'hEA8, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hFB9, 12'hFB9, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFB9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hEA8, 12'hE98, 12'hE97, 12'hE87, 12'hD87, 12'hD86, 12'hD76, 12'hC76, 12'hC87, 12'hE98, 12'hD88, 12'hE98, 12'hF98, 12'hFA8, 12'hFB9, 12'hFB9, 12'hFBA, 12'hFCB, 12'hFDB, 12'hFDC, 12'hFCB, 12'hFCB, 12'hFCB, 12'hFBA, 12'hFB9, 12'hFA9, 12'hFA8, 12'hE98, 12'hD87, 12'hC76, 12'hB65, 12'hA65, 12'h954, 12'h854, 12'h744, 12'h643, 12'h533, 12'h744, 12'h854, 12'h854, 12'h954, 12'h954, 12'h854, 12'h954, 12'h954, 12'h854, 12'h954, 12'h954, 12'h964, 12'h965, 12'h964, 12'h965, 12'h954, 12'h854, 12'h854, 12'h743, 12'h643, 12'h533, 12'h533, 12'h433, 12'h432, 12'h433, 12'h433, 12'h432, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h321, 12'h321, 12'h333, 12'hBBB, 12'hDDC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBC, 12'hCBB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBAB, 12'hBBA, 12'hBBB, 12'hBBB, 12'hBAA, 12'hABB, 12'hBBA,
		12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDDD, 12'hDBA, 12'hD98, 12'hD87, 12'hFBA, 12'hFA9, 12'hD86, 12'hC75, 12'hB64, 12'hB65, 12'hC75, 12'hD98, 12'hEAA, 12'hC98, 12'hC98, 12'hC97, 12'hC98, 12'hC98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hE98, 12'hEA8, 12'hD98, 12'hD98, 12'hEA8, 12'hEA8, 12'hEA9, 12'hEA9, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFB9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFB9, 12'hFA9, 12'hFA9, 12'hEA8, 12'hE97, 12'hE97, 12'hD87, 12'hD86, 12'hC76, 12'hC75, 12'hC76, 12'hD99, 12'hD88, 12'hE98, 12'hFA8, 12'hFB9, 12'hFCA, 12'hFDB, 12'hFDC, 12'hFDB, 12'hFDC, 12'hFDC, 12'hFED, 12'hFED, 12'hFED, 12'hFDC, 12'hFCB, 12'hFB9, 12'hFA8, 12'hFA8, 12'hFA8, 12'hD87, 12'hC76, 12'hB65, 12'hA65, 12'h954, 12'h854, 12'h854, 12'h754, 12'h643, 12'h643, 12'h855, 12'h865, 12'h965, 12'h954, 12'h854, 12'h954, 12'h954, 12'h954, 12'h964, 12'h954, 12'h954, 12'hA65, 12'h954, 12'hA65, 12'h954, 12'h954, 12'h854, 12'h754, 12'h643, 12'h643, 12'h543, 12'h433, 12'h433, 12'h432, 12'h433, 12'h432, 12'h333, 12'h333, 12'h332, 12'h322, 12'h322, 12'h322, 12'h321, 12'h322, 12'h989, 12'hDDD, 12'hDCD, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDC, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCDC, 12'hDCC, 12'hDBB, 12'hE99, 12'hC87, 12'hE97, 12'hFBA, 12'hF98, 12'hD86, 12'hB64, 12'hB64, 12'hB65, 12'hD87, 12'hDA9, 12'hC98, 12'hC87, 12'hD98, 12'hD98, 12'hC87, 12'hC87, 12'hC88, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD98, 12'hD97, 12'hE98, 12'hD97, 12'hE98, 12'hE98, 12'hE98, 12'hFA9, 12'hFA9, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFBA, 12'hFA9, 12'hFBA, 12'hFA9, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hEA8, 12'hE98, 12'hE97, 12'hE97, 12'hD87, 12'hD86, 12'hC76, 12'hC75, 12'hB76, 12'hC77, 12'hE99, 12'hE97, 12'hFA9, 12'hFB9, 12'hFCA, 12'hFCA, 12'hFBA, 12'hFA9, 12'hFA8, 12'hFA9, 12'hFB9, 12'hFBA, 12'hFCB, 12'hFCB, 12'hFCA, 12'hFB9, 12'hF98, 12'hF98, 12'hE97, 12'hE97, 12'hD86, 12'hB75, 12'h965, 12'h854, 12'h744, 12'h744, 12'h743, 12'h743, 12'h643, 12'h543, 12'h643, 12'h855, 12'h865, 12'h854, 12'h954, 12'h854, 12'h954, 12'h954, 12'h954, 12'h964, 12'h954, 12'h954, 12'h954, 12'h964, 12'h954, 12'h854, 12'h854, 12'h754, 12'h744, 12'h643, 12'h533, 12'h533, 12'h433, 12'h433, 12'h432, 12'h433, 12'h333, 12'h332, 12'h332, 12'h322, 12'h322, 12'h332, 12'h322, 12'h777, 12'hDDC, 12'hCCC, 12'hDDC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCBC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBA,
		12'hBCB, 12'hCCC, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hDCC, 12'hCDD, 12'hDDC, 12'hDDD, 12'hCDD, 12'hCDD, 12'hCCC, 12'hCCC, 12'hEA9, 12'hD87, 12'hC76, 12'hE98, 12'hFBA, 12'hFA8, 12'hE97, 12'hD75, 12'hB65, 12'hC87, 12'hC99, 12'hC98, 12'hC88, 12'hD98, 12'hD98, 12'hC87, 12'hC87, 12'hC98, 12'hC87, 12'hC87, 12'hD98, 12'hD98, 12'hD98, 12'hD87, 12'hC87, 12'hD97, 12'hD87, 12'hD98, 12'hE98, 12'hE98, 12'hEA8, 12'hFA9, 12'hFB9, 12'hFB9, 12'hFA9, 12'hFBA, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hEA8, 12'hFA9, 12'hE98, 12'hE98, 12'hD97, 12'hE87, 12'hD76, 12'hC76, 12'hC76, 12'hB65, 12'hC76, 12'hC88, 12'hD98, 12'hE97, 12'hFA8, 12'hFA8, 12'hF97, 12'hE76, 12'hA54, 12'h522, 12'h421, 12'h632, 12'hB65, 12'hF97, 12'hFA8, 12'hFA8, 12'hFA8, 12'hF97, 12'hF87, 12'hE76, 12'hD87, 12'hC86, 12'hB65, 12'h854, 12'h633, 12'h532, 12'h432, 12'h321, 12'h422, 12'h532, 12'h533, 12'h533, 12'h533, 12'h744, 12'h854, 12'h855, 12'h854, 12'h854, 12'h955, 12'h964, 12'h954, 12'h954, 12'h954, 12'h854, 12'h954, 12'h965, 12'h954, 12'h854, 12'h854, 12'h743, 12'h743, 12'h643, 12'h433, 12'h533, 12'h433, 12'h433, 12'h433, 12'h333, 12'h433, 12'h322, 12'h332, 12'h322, 12'h322, 12'h332, 12'h333, 12'hCCC, 12'hDDD, 12'hCDC, 12'hDCC, 12'hDCD, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCBB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hBCC, 12'hBCB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hDCD, 12'hDDC, 12'hCDC, 12'hCCC, 12'hDAA, 12'hE98, 12'hD86, 12'hD86, 12'hFA8, 12'hFBA, 12'hFB9, 12'hFA9, 12'hEBA, 12'hFDB, 12'hC98, 12'hC98, 12'hD98, 12'hC98, 12'hC87, 12'hC98, 12'hB87, 12'hB87, 12'hC98, 12'hC87, 12'hD98, 12'hB87, 12'hD87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hD97, 12'hD98, 12'hD97, 12'hEA8, 12'hEA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA8, 12'hFA9, 12'hFA8, 12'hFA8, 12'hEA8, 12'hE98, 12'hE98, 12'hE87, 12'hD87, 12'hD86, 12'hD76, 12'hC76, 12'hC75, 12'hC76, 12'hC76, 12'hD87, 12'hD99, 12'hD98, 12'hE88, 12'hE97, 12'hE87, 12'hC76, 12'h843, 12'h310, 12'h210, 12'h211, 12'h211, 12'h311, 12'h633, 12'hB66, 12'hF98, 12'hF97, 12'hF86, 12'hC65, 12'hB65, 12'hB66, 12'hA65, 12'h854, 12'h533, 12'h321, 12'h110, 12'h100, 12'h000, 12'h110, 12'h321, 12'h432, 12'h432, 12'h422, 12'h643, 12'h754, 12'h855, 12'h855, 12'h965, 12'h854, 12'h854, 12'h954, 12'h954, 12'h854, 12'h954, 12'h854, 12'h954, 12'h854, 12'h854, 12'h743, 12'h743, 12'h643, 12'h643, 12'h543, 12'h433, 12'h433, 12'h432, 12'h433, 12'h433, 12'h333, 12'h332, 12'h322, 12'h332, 12'h322, 12'h322, 12'h555, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDD, 12'hCDC, 12'hDDC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hBBC, 12'hCBB, 12'hCBB, 12'hBBB, 12'hCCB, 12'hCBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDCC, 12'hCDC, 12'hCCD, 12'hCCC, 12'hDCC, 12'hCDC, 12'hCCC, 12'hDBB, 12'hEB9, 12'hE98, 12'hD87, 12'hE87, 12'hF98, 12'hFA9, 12'hFBA, 12'hFCA, 12'hFBA, 12'hC87, 12'hC98, 12'hC98, 12'hC87, 12'hB87, 12'hC98, 12'hC98, 12'hC87, 12'hC87, 12'hC88, 12'hC87, 12'hC87, 12'hB86, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hC86, 12'hC77, 12'hD87, 12'hE98, 12'hE98, 12'hFA8, 12'hEA9, 12'hEA8, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFA8, 12'hFA8, 12'hE98, 12'hE98, 12'hE97, 12'hD87, 12'hD86, 12'hD86, 12'hC76, 12'hC76, 12'hC75, 12'hC76, 12'hC76, 12'hD88, 12'hD98, 12'hEA9, 12'hD99, 12'hD87, 12'hD87, 12'hC76, 12'hA54, 12'h632, 12'h421, 12'h421, 12'h422, 12'h422, 12'h633, 12'hA77, 12'hA77, 12'hA65, 12'hC76, 12'hB65, 12'h954, 12'h854, 12'h854, 12'h854, 12'h432, 12'h111, 12'h100, 12'h001, 12'h101, 12'h110, 12'h210, 12'h311, 12'h321, 12'h321, 12'h321, 12'h432, 12'h644, 12'h744, 12'h854, 12'h754, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h854, 12'h743, 12'h743, 12'h644, 12'h643, 12'h543, 12'h543, 12'h433, 12'h433, 12'h333, 12'h433, 12'h432, 12'h333, 12'h333, 12'h332, 12'h322, 12'h332, 12'h322, 12'h888, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDCD, 12'hDDD, 12'hDDD, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCBB, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCCC, 12'hBCB, 12'hBBB, 12'hCCC, 12'hCCB, 12'hBCC, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hCCC, 12'hCCC, 12'hBBB, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDBA, 12'hFA9, 12'hE97, 12'hD87, 12'hE98, 12'hFBA, 12'hFDB, 12'hFBA, 12'hFBA, 12'hC87, 12'hC98, 12'hD98, 12'hC98, 12'hC88, 12'hC98, 12'hC98, 12'hC98, 12'hC87, 12'hC87, 12'hB87, 12'hB87, 12'hB76, 12'hC87, 12'hB87, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hD87, 12'hD97, 12'hE98, 12'hE98, 12'hEA8, 12'hE98, 12'hE99, 12'hEA9, 12'hE98, 12'hE98, 12'hE98, 12'hE97, 12'hD86, 12'hD86, 12'hC76, 12'hC76, 12'hC76, 12'hB75, 12'hC76, 12'hC76, 12'hD88, 12'hE98, 12'hEA9, 12'hEAA, 12'hEAA, 12'hD99, 12'hC77, 12'hB65, 12'h954, 12'h844, 12'h844, 12'h965, 12'hC88, 12'hD98, 12'hD98, 12'hC88, 12'hB76, 12'hB76, 12'hB76, 12'h955, 12'h743, 12'h643, 12'h643, 12'h322, 12'h110, 12'h100, 12'h110, 12'h110, 12'h110, 12'h211, 12'h322, 12'h322, 12'h321, 12'h210, 12'h210, 12'h422, 12'h643, 12'h744, 12'h744, 12'h854, 12'h844, 12'h744, 12'h754, 12'h854, 12'h844, 12'h854, 12'h854, 12'h743, 12'h744, 12'h743, 12'h743, 12'h644, 12'h643, 12'h543, 12'h433, 12'h433, 12'h332, 12'h332, 12'h433, 12'h332, 12'h333, 12'h322, 12'h322, 12'h333, 12'h322, 12'h322, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDCD, 12'hDDC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCBC, 12'hCBB, 12'hCBC, 12'hCBB, 12'hCBB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCBC, 12'hCCC, 12'hCCB, 12'hCCB, 12'hBCC,
		12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCB, 12'hFAA, 12'hFA9, 12'hE97, 12'hEA9, 12'hFCA, 12'hFA8, 12'hE98, 12'hD98, 12'hC87, 12'hC98, 12'hB87, 12'hC98, 12'hC87, 12'hC87, 12'hC87, 12'hC98, 12'hC87, 12'hB77, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hA76, 12'hA65, 12'hA76, 12'hB76, 12'hC86, 12'hD87, 12'hD97, 12'hEA8, 12'hE98, 12'hE98, 12'hE98, 12'hEA8, 12'hE98, 12'hD98, 12'hD97, 12'hD87, 12'hC86, 12'hC76, 12'hB65, 12'hB75, 12'hB65, 12'hB65, 12'hB76, 12'hC87, 12'hE99, 12'hEA9, 12'hFA9, 12'hFBA, 12'hFA9, 12'hFA9, 12'hEA9, 12'hD99, 12'hC87, 12'hB77, 12'hD99, 12'hEA9, 12'hEAA, 12'hEAA, 12'hD98, 12'hD98, 12'hD98, 12'hC87, 12'hB77, 12'hA66, 12'h644, 12'h533, 12'h321, 12'h210, 12'h210, 12'h211, 12'h210, 12'h210, 12'h210, 12'h211, 12'h321, 12'h321, 12'h210, 12'h210, 12'h321, 12'h432, 12'h533, 12'h743, 12'h744, 12'h854, 12'h854, 12'h844, 12'h854, 12'h854, 12'h743, 12'h854, 12'h853, 12'h854, 12'h743, 12'h643, 12'h643, 12'h643, 12'h543, 12'h433, 12'h433, 12'h433, 12'h332, 12'h332, 12'h333, 12'h433, 12'h332, 12'h322, 12'h333, 12'h332, 12'h322, 12'h666, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCBC, 12'hCCB, 12'hCBC, 12'hBBB, 12'hCCB, 12'hCCC, 12'hBBB, 12'hCCC, 12'hBCB, 12'hBBB,
		12'hCCC, 12'hCCB, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDBA, 12'hFA9, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFA8, 12'hD98, 12'hEAA, 12'hB87, 12'hB88, 12'hB87, 12'hC87, 12'hC98, 12'hC87, 12'hC98, 12'hD98, 12'hC87, 12'hB87, 12'hA76, 12'hB76, 12'hB76, 12'hA76, 12'hB76, 12'hB76, 12'hA65, 12'hA76, 12'h965, 12'hB76, 12'hC86, 12'hC87, 12'hC87, 12'hD88, 12'hD98, 12'hD98, 12'hE98, 12'hD87, 12'hD98, 12'hD87, 12'hC87, 12'hC77, 12'hC76, 12'hB65, 12'hA65, 12'hA65, 12'hA66, 12'hB76, 12'hC87, 12'hD98, 12'hE99, 12'hEA9, 12'hFA9, 12'hFBA, 12'hFAA, 12'hFA9, 12'hFB9, 12'hFA9, 12'hFAA, 12'hFA9, 12'hEA9, 12'hFA9, 12'hFAA, 12'hEA9, 12'hDA9, 12'hD98, 12'hD88, 12'hC87, 12'hC87, 12'hB76, 12'h965, 12'h744, 12'h633, 12'h432, 12'h322, 12'h422, 12'h321, 12'h322, 12'h321, 12'h321, 12'h321, 12'h321, 12'h422, 12'h432, 12'h532, 12'h532, 12'h533, 12'h643, 12'h643, 12'h743, 12'h854, 12'h854, 12'h854, 12'h743, 12'h743, 12'h744, 12'h743, 12'h743, 12'h643, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h433, 12'h432, 12'h333, 12'h433, 12'h433, 12'h333, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCB, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBCC, 12'hBCB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hDDC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCDC, 12'hCDC, 12'hDBA, 12'hFBB, 12'hFA9, 12'hEA8, 12'hE99, 12'hEBA, 12'hFBA, 12'hC88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hC87, 12'hC87, 12'hC98, 12'hC87, 12'hB87, 12'hB76, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'hA66, 12'h965, 12'h965, 12'h965, 12'hB76, 12'hB76, 12'hB77, 12'hC87, 12'hD97, 12'hD98, 12'hD87, 12'hD88, 12'hC87, 12'hB77, 12'hB76, 12'hA65, 12'hA66, 12'hA66, 12'hA66, 12'hB76, 12'hB76, 12'hC87, 12'hD88, 12'hD98, 12'hE99, 12'hEA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hFA9, 12'hEA9, 12'hEA9, 12'hE99, 12'hEA9, 12'hDA9, 12'hD99, 12'hC98, 12'hC98, 12'hB87, 12'hC87, 12'hC87, 12'hC98, 12'hB87, 12'h966, 12'h855, 12'h644, 12'h644, 12'h644, 12'h433, 12'h533, 12'h532, 12'h633, 12'h633, 12'h633, 12'h633, 12'h643, 12'h633, 12'h633, 12'h633, 12'h533, 12'h633, 12'h643, 12'h744, 12'h744, 12'h744, 12'h743, 12'h743, 12'h744, 12'h643, 12'h643, 12'h633, 12'h533, 12'h533, 12'h543, 12'h433, 12'h432, 12'h332, 12'h333, 12'h332, 12'h332, 12'h322, 12'h322, 12'h232, 12'h322, 12'h333, 12'h665, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDCC, 12'hCDC, 12'hDCD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCBC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCCB, 12'hCBC, 12'hBCC, 12'hCCB, 12'hCBC, 12'hCCB, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hDDC, 12'hDDD, 12'hCCD, 12'hDDC, 12'hCDC, 12'hCCC, 12'hDDC, 12'hCCC, 12'hDCC, 12'hDDC, 12'hDDD, 12'hDCB, 12'hFB9, 12'hFBA, 12'hFBA, 12'hFCC, 12'hFBA, 12'hEA9, 12'hB87, 12'hB97, 12'hB87, 12'hC88, 12'hA76, 12'hC87, 12'hC87, 12'hB87, 12'hC88, 12'hC87, 12'hB87, 12'hB77, 12'hB76, 12'h965, 12'h965, 12'hA76, 12'hA75, 12'h965, 12'h965, 12'h965, 12'hA66, 12'hA76, 12'hC87, 12'hC87, 12'hD98, 12'hD98, 12'hC87, 12'hC87, 12'hA76, 12'hA76, 12'hA66, 12'hA76, 12'hA65, 12'hA76, 12'hB77, 12'hC87, 12'hC87, 12'hD88, 12'hD98, 12'hD98, 12'hE98, 12'hEA9, 12'hFA9, 12'hFA9, 12'hEA9, 12'hFA9, 12'hEA9, 12'hEA9, 12'hD98, 12'hD98, 12'hC88, 12'hDA9, 12'hC98, 12'hD99, 12'hC98, 12'hC98, 12'hD98, 12'hC88, 12'hC88, 12'hB77, 12'hC87, 12'hA76, 12'hA76, 12'h865, 12'h754, 12'h644, 12'h754, 12'h754, 12'h533, 12'h533, 12'h543, 12'h643, 12'h643, 12'h633, 12'h643, 12'h643, 12'h643, 12'h642, 12'h643, 12'h633, 12'h533, 12'h643, 12'h643, 12'h744, 12'h743, 12'h643, 12'h643, 12'h633, 12'h533, 12'h533, 12'h543, 12'h433, 12'h433, 12'h332, 12'h332, 12'h333, 12'h332, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h232, 12'h322, 12'hBBB, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCBC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hBCC, 12'hCCB, 12'hBBC, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hBBB, 12'hBCB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hDCD, 12'hDDD, 12'hCDD, 12'hDDD, 12'hDCC, 12'hCCC, 12'hCDC, 12'hCCD, 12'hDCC, 12'hCDD, 12'hDCC, 12'hEA9, 12'hFBA, 12'hFBA, 12'hFB9, 12'hFA8, 12'hD86, 12'hB77, 12'hA77, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hC87, 12'hB87, 12'hB87, 12'hC87, 12'hC87, 12'hB86, 12'hB76, 12'h965, 12'h965, 12'hA76, 12'h965, 12'h965, 12'h855, 12'h855, 12'hA76, 12'hA76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hB77, 12'hA66, 12'hA66, 12'hA76, 12'hA66, 12'hA76, 12'hB87, 12'hB87, 12'hB87, 12'hC88, 12'hC88, 12'hD98, 12'hD98, 12'hEA9, 12'hE98, 12'hEA9, 12'hD98, 12'hDA9, 12'hD98, 12'hD98, 12'hC98, 12'hC98, 12'hC98, 12'hC99, 12'hDA9, 12'hC98, 12'hC98, 12'hC88, 12'hB87, 12'hB87, 12'hC87, 12'hB87, 12'hB87, 12'hA76, 12'hB77, 12'hA76, 12'h965, 12'h855, 12'h854, 12'h643, 12'h854, 12'h754, 12'h643, 12'h533, 12'h533, 12'h532, 12'h643, 12'h643, 12'h643, 12'h633, 12'h643, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h643, 12'h643, 12'h643, 12'h533, 12'h533, 12'h533, 12'h433, 12'h433, 12'h432, 12'h432, 12'h332, 12'h332, 12'h323, 12'h322, 12'h332, 12'h323, 12'h332, 12'h222, 12'h222, 12'h222, 12'h444, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCD, 12'hCDC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCB, 12'hCCC, 12'hCBB, 12'hCCB, 12'hBBB, 12'hCBB, 12'hCCC, 12'hBBB, 12'hCCC, 12'hCCB, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hCBC, 12'hCBB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hCDC, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCDC, 12'hCCC, 12'hDCD, 12'hCDC, 12'hCDD, 12'hDDC, 12'hDCC, 12'hCCD, 12'hDDD, 12'hCAA, 12'hD87, 12'hE97, 12'hE87, 12'hD86, 12'hB64, 12'hA76, 12'hA76, 12'hB77, 12'hA77, 12'hA76, 12'hA77, 12'hB87, 12'hC87, 12'hB77, 12'hC87, 12'hC87, 12'hB87, 12'hA65, 12'h965, 12'h855, 12'h965, 12'h965, 12'h955, 12'h854, 12'h754, 12'h965, 12'hB76, 12'hB76, 12'hB87, 12'hC87, 12'hC88, 12'hB87, 12'hA76, 12'hA76, 12'h976, 12'h966, 12'h967, 12'h977, 12'hA87, 12'hA77, 12'hA77, 12'hB88, 12'hB88, 12'hC98, 12'hC98, 12'hC98, 12'hD98, 12'hB87, 12'hC98, 12'hC98, 12'hD98, 12'hC98, 12'hC88, 12'hC99, 12'hC88, 12'hC99, 12'hD98, 12'hDA9, 12'hC98, 12'hD98, 12'hC98, 12'hB87, 12'hB87, 12'hA76, 12'hA76, 12'hB76, 12'hA76, 12'hA76, 12'hA66, 12'h854, 12'h754, 12'h754, 12'h744, 12'h753, 12'h643, 12'h533, 12'h533, 12'h432, 12'h432, 12'h643, 12'h643, 12'h633, 12'h543, 12'h533, 12'h533, 12'h543, 12'h633, 12'h643, 12'h533, 12'h543, 12'h533, 12'h533, 12'h433, 12'h432, 12'h432, 12'h433, 12'h332, 12'h432, 12'h322, 12'h332, 12'h332, 12'h333, 12'h322, 12'h332, 12'h322, 12'h322, 12'h222, 12'h332, 12'h888, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDCC, 12'hCCC, 12'hDCD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCBC, 12'hCBB, 12'hCCC, 12'hCBC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCC, 12'hBCB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hBCB, 12'hCCC, 12'hCBC, 12'hBCB, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDD, 12'hDCC, 12'hCDD, 12'hDDC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hDCD, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDDC, 12'hDCC, 12'hCA9, 12'hB98, 12'hA87, 12'h866, 12'h866, 12'h976, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'hB87, 12'hC76, 12'hB87, 12'hB87, 12'hC87, 12'hB76, 12'hA76, 12'h955, 12'h754, 12'h854, 12'h965, 12'hA65, 12'h855, 12'h744, 12'h755, 12'hA66, 12'hC87, 12'hC87, 12'hC87, 12'hB77, 12'hB77, 12'hB87, 12'hA76, 12'hA76, 12'h967, 12'hA87, 12'hA77, 12'hA77, 12'hA88, 12'hA77, 12'hA87, 12'hB87, 12'hB88, 12'hB88, 12'hB88, 12'hC98, 12'hB88, 12'hD98, 12'hEA9, 12'hD99, 12'hC98, 12'hB88, 12'hB87, 12'hC98, 12'hC98, 12'hC88, 12'hC98, 12'hC88, 12'hC98, 12'hC97, 12'hB87, 12'hB77, 12'hA76, 12'hB87, 12'hB76, 12'hB87, 12'h976, 12'h965, 12'h855, 12'h754, 12'h754, 12'h644, 12'h543, 12'h543, 12'h643, 12'h543, 12'h432, 12'h432, 12'h433, 12'h433, 12'h432, 12'h433, 12'h533, 12'h533, 12'h533, 12'h533, 12'h543, 12'h433, 12'h533, 12'h533, 12'h533, 12'h433, 12'h432, 12'h432, 12'h433, 12'h332, 12'h332, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h322, 12'h222, 12'h222, 12'h332, 12'h222, 12'hAAA, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDCD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCCC, 12'hBBB, 12'hCCB, 12'hCCC, 12'hBBB, 12'hCCB, 12'hBBC, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBBB, 12'hCCB, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDC, 12'hCCD, 12'hCDC, 12'hCCD, 12'hDCD, 12'hCDC, 12'hCDC, 12'hDCC, 12'hCCC, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hA99, 12'h988, 12'h966, 12'hA87, 12'h976, 12'hA66, 12'hA76, 12'hA76, 12'hB76, 12'hB76, 12'hB76, 12'hB76, 12'hC87, 12'hB76, 12'hA76, 12'h855, 12'h754, 12'h865, 12'h965, 12'hA65, 12'h754, 12'h755, 12'hA76, 12'hC87, 12'hC87, 12'hC88, 12'hB87, 12'hA77, 12'hB87, 12'h977, 12'hA77, 12'hA77, 12'hA77, 12'h977, 12'hA77, 12'hA87, 12'h977, 12'hA77, 12'hA87, 12'hB88, 12'hB87, 12'hC88, 12'hB88, 12'hC88, 12'hC98, 12'hC88, 12'hD98, 12'hC98, 12'hC98, 12'hD99, 12'hD98, 12'hDA9, 12'hEA9, 12'hEA9, 12'hEA9, 12'hE99, 12'hE98, 12'hD98, 12'hC87, 12'hB76, 12'hC87, 12'hB76, 12'hB87, 12'hB87, 12'hB76, 12'hB76, 12'h965, 12'h744, 12'h643, 12'h543, 12'h533, 12'h433, 12'h432, 12'h432, 12'h432, 12'h322, 12'h322, 12'h433, 12'h332, 12'h433, 12'h432, 12'h432, 12'h433, 12'h433, 12'h543, 12'h432, 12'h543, 12'h533, 12'h433, 12'h332, 12'h332, 12'h332, 12'h322, 12'h332, 12'h322, 12'h332, 12'h332, 12'h222, 12'h322, 12'h322, 12'h222, 12'h222, 12'h322, 12'h332, 12'h666, 12'hDDD, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCBC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCBC, 12'hBCB, 12'hBBB, 12'hBBC, 12'hCCB, 12'hBCB, 12'hBBC, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hBBC, 12'hBBB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCD, 12'hCDC, 12'hCCC, 12'hDDD, 12'hDCC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hDDC, 12'hDCC, 12'hCCC, 12'hCBB, 12'hBAA, 12'h766, 12'hA77, 12'hA77, 12'h966, 12'h966, 12'h965, 12'hA76, 12'hA76, 12'hB76, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hA76, 12'h965, 12'h855, 12'h755, 12'h966, 12'hA76, 12'h966, 12'h855, 12'hA76, 12'hC86, 12'hD98, 12'hB87, 12'hB88, 12'hB87, 12'hA77, 12'hA77, 12'h977, 12'h966, 12'h976, 12'h976, 12'h867, 12'h866, 12'h756, 12'h866, 12'h866, 12'hA77, 12'hA88, 12'hB88, 12'hC98, 12'hD98, 12'hD98, 12'hEA9, 12'hEA9, 12'hEA9, 12'hEBA, 12'hEAA, 12'hFA9, 12'hFAA, 12'hEA9, 12'hEA9, 12'hE99, 12'hE99, 12'hE99, 12'hE98, 12'hE98, 12'hD87, 12'hC87, 12'hD87, 12'hD87, 12'hC87, 12'hC86, 12'hC76, 12'hA65, 12'h965, 12'h854, 12'h744, 12'h643, 12'h533, 12'h322, 12'h422, 12'h322, 12'h322, 12'h322, 12'h321, 12'h322, 12'h322, 12'h222, 12'h322, 12'h332, 12'h432, 12'h433, 12'h332, 12'h433, 12'h543, 12'h433, 12'h322, 12'h332, 12'h433, 12'h322, 12'h322, 12'h332, 12'h322, 12'h322, 12'h332, 12'h222, 12'h332, 12'h322, 12'h222, 12'h222, 12'h332, 12'h545, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hCBB, 12'hBBB,
		12'hBBB, 12'hBCB, 12'hCBB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hDDD, 12'hDDC, 12'hCCC, 12'hDDD, 12'hDCC, 12'hDCC, 12'hDDD, 12'hCCC, 12'hBBB, 12'h988, 12'h888, 12'h877, 12'h977, 12'h865, 12'h965, 12'h976, 12'hA76, 12'hA76, 12'h966, 12'hB76, 12'hA76, 12'hC87, 12'hB86, 12'hC87, 12'hB87, 12'hB77, 12'hB76, 12'h966, 12'h965, 12'hA66, 12'hA77, 12'h976, 12'hA76, 12'hC87, 12'hC98, 12'hC88, 12'hC88, 12'hB87, 12'hB77, 12'hA77, 12'h966, 12'h966, 12'h966, 12'h866, 12'h755, 12'h655, 12'h655, 12'h866, 12'hA77, 12'hB88, 12'hC98, 12'hD98, 12'hEA9, 12'hEA9, 12'hD99, 12'hE99, 12'hD99, 12'hD99, 12'hD98, 12'hD88, 12'hC88, 12'hC88, 12'hC88, 12'hC87, 12'hC87, 12'hC88, 12'hC77, 12'hB77, 12'hB77, 12'hB67, 12'hB66, 12'hA65, 12'hA55, 12'h954, 12'h844, 12'h744, 12'h743, 12'h733, 12'h643, 12'h743, 12'h743, 12'h643, 12'h533, 12'h543, 12'h332, 12'h333, 12'h322, 12'h321, 12'h221, 12'h221, 12'h221, 12'h221, 12'h222, 12'h322, 12'h432, 12'h322, 12'h322, 12'h443, 12'h533, 12'h433, 12'h433, 12'h432, 12'h332, 12'h232, 12'h322, 12'h322, 12'h332, 12'h222, 12'h222, 12'h322, 12'h222, 12'h222, 12'h232, 12'h322, 12'h766, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCB, 12'hDCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBBB, 12'hCBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hCCB, 12'hBCB, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hDDD, 12'hDDD, 12'hDCD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCBB, 12'hCBB, 12'h988, 12'h777, 12'h555, 12'h977, 12'h966, 12'h976, 12'h865, 12'h966, 12'hA77, 12'h966, 12'hA76, 12'h965, 12'hB76, 12'hB76, 12'hA76, 12'hC87, 12'hC87, 12'hA76, 12'hA77, 12'h966, 12'hB76, 12'hA77, 12'h977, 12'hA76, 12'hB76, 12'hD88, 12'hC87, 12'hC87, 12'hC88, 12'hA87, 12'hA77, 12'h966, 12'h866, 12'h866, 12'h755, 12'h755, 12'h644, 12'h654, 12'h755, 12'h655, 12'h633, 12'h744, 12'h955, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hB67, 12'hB77, 12'hB77, 12'hC88, 12'hB77, 12'hB77, 12'hC78, 12'hC88, 12'hC78, 12'hB77, 12'hB88, 12'hB77, 12'hB77, 12'hA77, 12'hA66, 12'h855, 12'h745, 12'h755, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h422, 12'h422, 12'h432, 12'h422, 12'h322, 12'h422, 12'h322, 12'h321, 12'h221, 12'h211, 12'h111, 12'h111, 12'h211, 12'h222, 12'h222, 12'h332, 12'h322, 12'h333, 12'h533, 12'h433, 12'h433, 12'h432, 12'h332, 12'h322, 12'h222, 12'h232, 12'h332, 12'h222, 12'h322, 12'h322, 12'h222, 12'h222, 12'h322, 12'h232, 12'h555, 12'hCCC, 12'hDDD, 12'hEED, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBCC, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hCBB, 12'hBCC, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCDC, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDCD, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hAAA, 12'h988, 12'h666, 12'h876, 12'h976, 12'h976, 12'h966, 12'h966, 12'h965, 12'h966, 12'h965, 12'h965, 12'hA76, 12'hA65, 12'hB76, 12'hB76, 12'hB87, 12'hC98, 12'hA77, 12'hA77, 12'hA77, 12'hB88, 12'h977, 12'hB77, 12'hB77, 12'hC87, 12'hC88, 12'hC88, 12'hC88, 12'hB87, 12'hA77, 12'h966, 12'h865, 12'h866, 12'h755, 12'h765, 12'h765, 12'h856, 12'h977, 12'hA77, 12'hB88, 12'h855, 12'h966, 12'h956, 12'h845, 12'h855, 12'h855, 12'h966, 12'h855, 12'h956, 12'h966, 12'h966, 12'h966, 12'h966, 12'h966, 12'hA66, 12'h966, 12'hA77, 12'hA66, 12'hA66, 12'hA66, 12'h955, 12'h744, 12'h744, 12'h643, 12'h533, 12'h533, 12'h422, 12'h322, 12'h322, 12'h322, 12'h222, 12'h211, 12'h211, 12'h211, 12'h210, 12'h210, 12'h111, 12'h110, 12'h111, 12'h211, 12'h211, 12'h222, 12'h322, 12'h322, 12'h433, 12'h433, 12'h433, 12'h443, 12'h433, 12'h433, 12'h332, 12'h333, 12'h322, 12'h322, 12'h333, 12'h332, 12'h322, 12'h222, 12'h322, 12'h222, 12'h222, 12'h222, 12'h666, 12'hEEE, 12'hDDD, 12'hEDD, 12'hEEE, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCBC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hCCC, 12'hBBB, 12'hCBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hCCB, 12'hCBC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hDDC, 12'hDDD, 12'hCDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCD, 12'hDCC, 12'hCCC, 12'hCBB, 12'hBAA, 12'h666, 12'h866, 12'hA77, 12'h966, 12'h977, 12'h866, 12'h976, 12'h965, 12'h965, 12'h966, 12'h965, 12'hA65, 12'hB76, 12'hC87, 12'hC87, 12'hC88, 12'hC98, 12'hB88, 12'hA77, 12'hB88, 12'hA77, 12'h966, 12'hB87, 12'hC88, 12'hC88, 12'hC98, 12'hC88, 12'hB87, 12'h977, 12'h977, 12'h755, 12'h866, 12'h755, 12'h866, 12'h866, 12'h866, 12'h966, 12'hA77, 12'hC88, 12'hD99, 12'hC88, 12'hC78, 12'hC78, 12'hC77, 12'hC67, 12'hB56, 12'h945, 12'h844, 12'h533, 12'h533, 12'h634, 12'h634, 12'h856, 12'h855, 12'h855, 12'h845, 12'h855, 12'h745, 12'h744, 12'h744, 12'h533, 12'h533, 12'h533, 12'h422, 12'h322, 12'h321, 12'h211, 12'h210, 12'h211, 12'h210, 12'h211, 12'h210, 12'h110, 12'h110, 12'h110, 12'h111, 12'h221, 12'h322, 12'h222, 12'h322, 12'h332, 12'h332, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h332, 12'h332, 12'h333, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h221, 12'h332, 12'hBBB, 12'hDDD, 12'hEDD, 12'hDEE, 12'hEDE, 12'hDDD, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCCC, 12'hBCB, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBBC, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hCCC, 12'hCBB, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hDDD, 12'hCCD, 12'hDDC, 12'hDDC, 12'hCDD, 12'hDCC, 12'hDCC, 12'hCBB, 12'hCBB, 12'h988, 12'h776, 12'h755, 12'hA77, 12'h976, 12'h966, 12'h866, 12'h865, 12'h966, 12'h865, 12'h965, 12'h966, 12'h965, 12'hA76, 12'hB77, 12'hB76, 12'hB87, 12'hB77, 12'hB88, 12'hB87, 12'hC98, 12'hA88, 12'h966, 12'hA77, 12'hB87, 12'hC87, 12'hC98, 12'hB77, 12'hA77, 12'hA77, 12'hA76, 12'h755, 12'h756, 12'h866, 12'h866, 12'h866, 12'h966, 12'hA77, 12'hA77, 12'hC88, 12'hD98, 12'hD99, 12'hEAA, 12'hD9A, 12'hD78, 12'hD89, 12'hE89, 12'hE89, 12'hD78, 12'hD78, 12'hC67, 12'hA56, 12'hB67, 12'hC78, 12'hC67, 12'hB67, 12'hA56, 12'h955, 12'h845, 12'h844, 12'h734, 12'h623, 12'h633, 12'h633, 12'h633, 12'h523, 12'h523, 12'h533, 12'h533, 12'h422, 12'h422, 12'h422, 12'h322, 12'h322, 12'h322, 12'h432, 12'h433, 12'h432, 12'h322, 12'h322, 12'h332, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h332, 12'h332, 12'h322, 12'h332, 12'h322, 12'h322, 12'h222, 12'h322, 12'h221, 12'h221, 12'h222, 12'h555, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDE, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCBB, 12'hCBB, 12'hBCC, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCB, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hCCC, 12'hCCC, 12'hDDD, 12'hCCC, 12'hDDC, 12'hDDD, 12'hCCC, 12'hBBB, 12'hA99, 12'h777, 12'h977, 12'hA77, 12'hA87, 12'h866, 12'h966, 12'h866, 12'h865, 12'h855, 12'h965, 12'h965, 12'h966, 12'hA75, 12'hB76, 12'hC86, 12'hC87, 12'hB87, 12'hB88, 12'hB88, 12'hC88, 12'hA88, 12'hA77, 12'hB87, 12'hB87, 12'hB87, 12'hB77, 12'hB87, 12'hB88, 12'hA76, 12'h866, 12'h866, 12'h866, 12'h966, 12'h866, 12'h966, 12'hA77, 12'hA77, 12'hA77, 12'hB77, 12'hC88, 12'hD98, 12'hD99, 12'hE9A, 12'hEAA, 12'hEAB, 12'hEAB, 12'hFAB, 12'hE9A, 12'hE9A, 12'hE89, 12'hE89, 12'hE89, 12'hE89, 12'hE89, 12'hE89, 12'hD78, 12'hD78, 12'hD78, 12'hD88, 12'hC77, 12'hB67, 12'hC78, 12'hC68, 12'hB67, 12'hA66, 12'hA56, 12'h955, 12'h955, 12'h745, 12'h644, 12'h634, 12'h534, 12'h544, 12'h433, 12'h433, 12'h422, 12'h322, 12'h322, 12'h322, 12'h322, 12'h433, 12'h333, 12'h433, 12'h433, 12'h443, 12'h444, 12'h443, 12'h333, 12'h433, 12'h332, 12'h333, 12'h322, 12'h222, 12'h332, 12'h222, 12'h322, 12'h221, 12'h322, 12'h222, 12'h222, 12'hBBB, 12'hDEE, 12'hDDD, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCCC, 12'hCBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB,
		12'hCBB, 12'hBCB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hBCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCBB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hCCC, 12'hCDD, 12'hCCC, 12'hDDD, 12'hCCC, 12'hCDD, 12'hDDD, 12'hCCC, 12'hBBB, 12'h988, 12'hB98, 12'hC98, 12'hA77, 12'h976, 12'h966, 12'h865, 12'h866, 12'h855, 12'h865, 12'h855, 12'hA66, 12'hA76, 12'hA65, 12'hB76, 12'hC87, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'hA77, 12'hA88, 12'hB87, 12'hB77, 12'hB77, 12'hA77, 12'h977, 12'hA77, 12'h966, 12'h866, 12'h866, 12'h866, 12'h966, 12'h977, 12'h977, 12'hA76, 12'hA77, 12'hB87, 12'hB77, 12'hA77, 12'hC88, 12'hC88, 12'hD98, 12'hE98, 12'hE99, 12'hEAB, 12'hFCC, 12'hFBC, 12'hFBC, 12'hFBC, 12'hFBC, 12'hFBB, 12'hFAB, 12'hFAB, 12'hF9A, 12'hE9A, 12'hE89, 12'hE8A, 12'hE89, 12'hD88, 12'hC67, 12'hD89, 12'hD78, 12'hC67, 12'hB67, 12'hB66, 12'hA56, 12'h945, 12'h845, 12'h744, 12'h644, 12'h533, 12'h533, 12'h432, 12'h322, 12'h322, 12'h322, 12'h432, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h433, 12'h433, 12'h433, 12'h332, 12'h332, 12'h222, 12'h332, 12'h322, 12'h222, 12'h222, 12'h221, 12'h221, 12'h222, 12'h555, 12'hEEE, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCB, 12'hCBC, 12'hCBB, 12'hCCB, 12'hBBB, 12'hCBB, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDDC, 12'hDDD, 12'hCCC, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCCB, 12'hA99, 12'hB98, 12'hDA9, 12'hA77, 12'h966, 12'h866, 12'h866, 12'h865, 12'h865, 12'h976, 12'h865, 12'h965, 12'h965, 12'hA76, 12'hB76, 12'hA66, 12'hA76, 12'hB77, 12'hA77, 12'hA87, 12'hA77, 12'hA77, 12'hA77, 12'hB87, 12'hA77, 12'h967, 12'h977, 12'hA76, 12'hA77, 12'h966, 12'h855, 12'h866, 12'h976, 12'h966, 12'h977, 12'hA77, 12'hA77, 12'hA87, 12'hB77, 12'hB77, 12'hA77, 12'hB77, 12'hC87, 12'hC88, 12'hD88, 12'hD88, 12'hD88, 12'hE99, 12'hE9A, 12'hFAB, 12'hFBC, 12'hFBC, 12'hFAB, 12'hEAB, 12'hFAB, 12'hEAA, 12'hE99, 12'hE89, 12'hE89, 12'hD89, 12'hC78, 12'hD88, 12'hC77, 12'hB66, 12'hB66, 12'hA56, 12'h955, 12'h845, 12'h744, 12'h644, 12'h533, 12'h432, 12'h422, 12'h322, 12'h322, 12'h322, 12'h332, 12'h433, 12'h433, 12'h433, 12'h443, 12'h433, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h322, 12'h222, 12'h322, 12'h221, 12'h221, 12'h222, 12'hAAA, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBCC, 12'hCBC, 12'hCCB, 12'hBBC, 12'hCBB, 12'hBBB, 12'hBCC, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hBBB, 12'hBCC, 12'hBCB, 12'hCBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hDDC, 12'hCCC, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBAA, 12'hCA9, 12'hDA9, 12'hB87, 12'hA77, 12'h966, 12'h976, 12'h866, 12'h866, 12'h855, 12'h965, 12'h965, 12'h965, 12'hA66, 12'h965, 12'hA66, 12'hA76, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'h966, 12'hB87, 12'hB77, 12'h977, 12'hA77, 12'h966, 12'h966, 12'h865, 12'h866, 12'h766, 12'h866, 12'h977, 12'hA78, 12'hB87, 12'hA77, 12'hB88, 12'hC88, 12'hC87, 12'hC98, 12'hB87, 12'hB77, 12'hC87, 12'hB87, 12'hB87, 12'hC87, 12'hC87, 12'hC77, 12'hC77, 12'hD77, 12'hD78, 12'hD88, 12'hD88, 12'hD89, 12'hD88, 12'hC78, 12'hD78, 12'hC78, 12'hB77, 12'hB67, 12'hB67, 12'hA66, 12'hA55, 12'h955, 12'h845, 12'h744, 12'h744, 12'h633, 12'h432, 12'h422, 12'h321, 12'h321, 12'h322, 12'h322, 12'h332, 12'h432, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h332, 12'h322, 12'h332, 12'h222, 12'h222, 12'h222, 12'h221, 12'h221, 12'h221, 12'h222, 12'h555, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDCC, 12'hDCD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCCC, 12'hBBB, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCBC, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDCC, 12'hCDC, 12'hDDD, 12'hCCC, 12'hDCC, 12'hCCC, 12'hBBB, 12'hBBB, 12'hDDD, 12'hDDD, 12'hDDC, 12'hBBB, 12'hCBB, 12'hDAA, 12'hDA9, 12'hD98, 12'h966, 12'h976, 12'hA77, 12'h966, 12'h966, 12'h866, 12'h855, 12'h855, 12'hA76, 12'h965, 12'hA76, 12'hA65, 12'hB76, 12'h965, 12'h966, 12'h966, 12'h977, 12'h976, 12'hA77, 12'hA76, 12'hA77, 12'h976, 12'h977, 12'h977, 12'h866, 12'h865, 12'h866, 12'h766, 12'h866, 12'h967, 12'h977, 12'hB88, 12'hA77, 12'h977, 12'hA77, 12'hB77, 12'hB87, 12'hB77, 12'hB77, 12'hB77, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'hA76, 12'hA66, 12'hA76, 12'hA65, 12'hA66, 12'hA66, 12'hA65, 12'h955, 12'h965, 12'h854, 12'h844, 12'h744, 12'h744, 12'h744, 12'h633, 12'h633, 12'h533, 12'h432, 12'h322, 12'h321, 12'h221, 12'h211, 12'h222, 12'h321, 12'h332, 12'h432, 12'h432, 12'h432, 12'h433, 12'h433, 12'h443, 12'h433, 12'h433, 12'h433, 12'h333, 12'h443, 12'h433, 12'h333, 12'h332, 12'h222, 12'h222, 12'h222, 12'h322, 12'h221, 12'h221, 12'h222, 12'h222, 12'h333, 12'hCCC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCCC, 12'hCBB, 12'hBCB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBCB, 12'hBCB, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBBB, 12'h989, 12'h888, 12'h888, 12'h777, 12'h666, 12'h888, 12'hA9A, 12'hBA9, 12'hDBA, 12'hDA9, 12'hEA9, 12'hA76, 12'h976, 12'h966, 12'h966, 12'h966, 12'h866, 12'h866, 12'h866, 12'h965, 12'h965, 12'hA66, 12'hA76, 12'hA66, 12'h976, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'hA77, 12'h966, 12'hA76, 12'hB77, 12'h966, 12'h645, 12'h866, 12'h866, 12'h755, 12'h867, 12'h877, 12'h867, 12'h977, 12'h977, 12'h976, 12'h976, 12'hA77, 12'hA77, 12'hB87, 12'hB77, 12'hC87, 12'hB87, 12'hB77, 12'hB77, 12'hB76, 12'hA76, 12'h866, 12'h855, 12'h655, 12'h755, 12'h754, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h755, 12'h543, 12'h533, 12'h332, 12'h322, 12'h332, 12'h322, 12'h322, 12'h322, 12'h221, 12'h211, 12'h222, 12'h221, 12'h321, 12'h322, 12'h322, 12'h432, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h544, 12'h444, 12'h443, 12'h444, 12'h333, 12'h443, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h211, 12'h222, 12'h222, 12'hAAB, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hCCD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBC, 12'hBCC, 12'hCCB, 12'hCCC, 12'hBBC, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBCB, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hBAB, 12'h989, 12'h888, 12'h989, 12'h888, 12'h666, 12'h434, 12'h656, 12'h878, 12'hBAA, 12'hDBA, 12'hD99, 12'hEA9, 12'hD98, 12'h976, 12'hA77, 12'h966, 12'hA76, 12'h966, 12'h966, 12'h865, 12'h755, 12'h865, 12'h965, 12'h965, 12'h966, 12'h865, 12'h966, 12'h966, 12'h966, 12'h965, 12'h966, 12'h966, 12'h966, 12'hA76, 12'hA66, 12'hA77, 12'h966, 12'h766, 12'h867, 12'h766, 12'h876, 12'hA77, 12'h977, 12'hA88, 12'h967, 12'h867, 12'h866, 12'hA87, 12'hB87, 12'hB87, 12'hB87, 12'hC87, 12'hB87, 12'hC87, 12'hB77, 12'hB77, 12'hA77, 12'hA76, 12'h966, 12'h855, 12'h865, 12'h755, 12'h755, 12'h654, 12'h544, 12'h544, 12'h644, 12'h544, 12'h433, 12'h423, 12'h433, 12'h433, 12'h332, 12'h322, 12'h321, 12'h322, 12'h322, 12'h321, 12'h322, 12'h422, 12'h432, 12'h432, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h443, 12'h433, 12'h443, 12'h433, 12'h433, 12'h433, 12'h433, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h221, 12'h111, 12'h222, 12'h222, 12'h999, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDCD, 12'hCCC, 12'hDDC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCB, 12'hBBB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hCBC, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hDDC, 12'hCCC, 12'hAAA, 12'h999, 12'h989, 12'h989, 12'h777, 12'h878, 12'h766, 12'h545, 12'h555, 12'h444, 12'hA88, 12'hDAA, 12'hDA9, 12'hD99, 12'hE98, 12'hB87, 12'h966, 12'h977, 12'h977, 12'h866, 12'h976, 12'h866, 12'h855, 12'h866, 12'h865, 12'h855, 12'h855, 12'h865, 12'h866, 12'h965, 12'h866, 12'h855, 12'h966, 12'h966, 12'h966, 12'hA76, 12'h966, 12'h966, 12'h866, 12'h866, 12'h866, 12'h866, 12'h867, 12'h866, 12'hA77, 12'h977, 12'h976, 12'h966, 12'h977, 12'hA77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB87, 12'hB77, 12'hC87, 12'hB77, 12'hB76, 12'hB76, 12'hA76, 12'h966, 12'h865, 12'h855, 12'h755, 12'h755, 12'h855, 12'h754, 12'h644, 12'h644, 12'h644, 12'h544, 12'h433, 12'h432, 12'h533, 12'h432, 12'h432, 12'h432, 12'h422, 12'h432, 12'h433, 12'h433, 12'h432, 12'h433, 12'h433, 12'h432, 12'h433, 12'h333, 12'h433, 12'h433, 12'h444, 12'h433, 12'h433, 12'h333, 12'h333, 12'h322, 12'h222, 12'h222, 12'h221, 12'h221, 12'h221, 12'h211, 12'h221, 12'h122, 12'h889, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDCD, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBBB, 12'hA9A, 12'h999, 12'h878, 12'h888, 12'h777, 12'h777, 12'h766, 12'h555, 12'h333, 12'h222, 12'h988, 12'hEBA, 12'hDA9, 12'hD98, 12'hE98, 12'hD98, 12'hA76, 12'h866, 12'h966, 12'h977, 12'h966, 12'h966, 12'h866, 12'h755, 12'h755, 12'h855, 12'h855, 12'h865, 12'h855, 12'h855, 12'h865, 12'h755, 12'h865, 12'h865, 12'h966, 12'h866, 12'h966, 12'h866, 12'h966, 12'h855, 12'h766, 12'h866, 12'h756, 12'h877, 12'h977, 12'h977, 12'h977, 12'hA87, 12'hA77, 12'hA77, 12'hA77, 12'hB87, 12'hB88, 12'hB77, 12'hB77, 12'hC87, 12'hC87, 12'hB77, 12'hB77, 12'hB76, 12'hB77, 12'hB77, 12'hB76, 12'hA66, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h754, 12'h754, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h432, 12'h533, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h332, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h332, 12'h322, 12'h222, 12'h222, 12'h221, 12'h221, 12'h211, 12'h111, 12'h221, 12'h222, 12'h989, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDC, 12'hCCD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hBCC, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBC, 12'hBBB, 12'hBCB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hCCC, 12'hCCB, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCDC, 12'hDCC, 12'hCBB, 12'h999, 12'hA9A, 12'h989, 12'h878, 12'h878, 12'h777, 12'h767, 12'h656, 12'h545, 12'h433, 12'h222, 12'h866, 12'hEBA, 12'hDA9, 12'hD98, 12'hDA9, 12'hEA8, 12'hC87, 12'h966, 12'h866, 12'h966, 12'h866, 12'h966, 12'h866, 12'h755, 12'h866, 12'h755, 12'h865, 12'h754, 12'h855, 12'h754, 12'h755, 12'h755, 12'h855, 12'h865, 12'h865, 12'h866, 12'h865, 12'h755, 12'h966, 12'h766, 12'h866, 12'h755, 12'h756, 12'h877, 12'h866, 12'hA88, 12'hA77, 12'h977, 12'hA87, 12'hA77, 12'hA88, 12'hB88, 12'hB87, 12'hB88, 12'hB88, 12'hB77, 12'hB87, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hB77, 12'hB76, 12'hA76, 12'h965, 12'h966, 12'h865, 12'h865, 12'h855, 12'h755, 12'h644, 12'h644, 12'h754, 12'h644, 12'h643, 12'h533, 12'h533, 12'h543, 12'h533, 12'h533, 12'h533, 12'h543, 12'h543, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h443, 12'h333, 12'h332, 12'h333, 12'h322, 12'h222, 12'h222, 12'h221, 12'h222, 12'h211, 12'h211, 12'h121, 12'h222, 12'h667, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hCCD, 12'hCCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hCCC, 12'hBCC, 12'hCCB, 12'hCCC, 12'hBCC, 12'hCDC, 12'hCDC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hCCC, 12'hCDC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hBBB, 12'hA9A, 12'h989, 12'hAAA, 12'h889, 12'h989, 12'hA99, 12'h878, 12'h767, 12'h766, 12'h666, 12'h434, 12'h111, 12'h766, 12'hDA9, 12'hEAA, 12'hD99, 12'hD98, 12'hD98, 12'hD98, 12'hB77, 12'h977, 12'h976, 12'h976, 12'h966, 12'h966, 12'h865, 12'h755, 12'h765, 12'h755, 12'h755, 12'h855, 12'h855, 12'h754, 12'h865, 12'h856, 12'h755, 12'h755, 12'h755, 12'h755, 12'h866, 12'h755, 12'h866, 12'h755, 12'h876, 12'h655, 12'h866, 12'h977, 12'h977, 12'h977, 12'hA77, 12'hB88, 12'h977, 12'hA88, 12'hA78, 12'hB88, 12'hC88, 12'hB88, 12'hB87, 12'hC88, 12'hC88, 12'hC88, 12'hC87, 12'hB87, 12'hB87, 12'hB76, 12'hB76, 12'hA77, 12'hA66, 12'hA76, 12'hA66, 12'hA66, 12'hA66, 12'h965, 12'h854, 12'h855, 12'h754, 12'h644, 12'h643, 12'h633, 12'h643, 12'h543, 12'h543, 12'h533, 12'h543, 12'h544, 12'h543, 12'h433, 12'h433, 12'h333, 12'h332, 12'h332, 12'h333, 12'h433, 12'h333, 12'h433, 12'h333, 12'h222, 12'h222, 12'h221, 12'h221, 12'h111, 12'h111, 12'h121, 12'h222, 12'h555, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDDC, 12'hDDC, 12'hDDD, 12'hCCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hBCC, 12'hCBC, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hCCC, 12'hBCB, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hDDC, 12'hCDC, 12'hCBC, 12'hBBB, 12'hA9A, 12'h99A, 12'hAAA, 12'h99A, 12'hAAA, 12'h999, 12'h888, 12'h999, 12'h888, 12'h989, 12'h767, 12'h878, 12'h877, 12'h555, 12'h322, 12'h644, 12'hCA9, 12'hDA9, 12'hD99, 12'hC88, 12'hD98, 12'hD98, 12'hD98, 12'hA77, 12'h866, 12'h977, 12'h966, 12'h966, 12'h766, 12'h855, 12'h755, 12'h755, 12'h755, 12'h754, 12'h754, 12'h755, 12'h644, 12'h755, 12'h544, 12'h644, 12'h755, 12'h755, 12'h654, 12'h755, 12'h755, 12'h866, 12'h866, 12'h866, 12'h977, 12'h977, 12'hA88, 12'h977, 12'hA78, 12'hB88, 12'hA88, 12'hC88, 12'hC88, 12'hB88, 12'hB87, 12'hB88, 12'hB77, 12'hC88, 12'hC87, 12'hC88, 12'hC88, 12'hC87, 12'hC87, 12'hC87, 12'hC87, 12'hB77, 12'hC87, 12'hB76, 12'hB76, 12'hB76, 12'hA66, 12'h955, 12'h865, 12'h855, 12'h754, 12'h643, 12'h643, 12'h644, 12'h533, 12'h644, 12'h644, 12'h643, 12'h644, 12'h544, 12'h533, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h332, 12'h332, 12'h333, 12'h433, 12'h322, 12'h222, 12'h222, 12'h221, 12'h111, 12'h121, 12'h111, 12'h222, 12'h777, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hBBC, 12'hBCB, 12'hBBB, 12'hCBB, 12'hBCC, 12'hBBB, 12'hBCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hBCB, 12'hBCB, 12'hCCC, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCD, 12'hCCD, 12'hBBB, 12'hA9A, 12'h878, 12'h878, 12'hAAA, 12'h989, 12'h989, 12'h99A, 12'h999, 12'h889, 12'h999, 12'h889, 12'h778, 12'h888, 12'h878, 12'h767, 12'h777, 12'h443, 12'h433, 12'hA88, 12'hD99, 12'hDA9, 12'hC87, 12'hC87, 12'hD98, 12'hD98, 12'hD97, 12'h976, 12'h967, 12'h976, 12'h977, 12'h866, 12'h866, 12'h866, 12'h855, 12'h654, 12'h654, 12'h754, 12'h654, 12'h655, 12'h654, 12'h755, 12'h655, 12'h644, 12'h644, 12'h755, 12'h644, 12'h655, 12'h755, 12'h755, 12'h866, 12'h866, 12'h977, 12'h977, 12'hA88, 12'hC98, 12'hC98, 12'hB88, 12'hC98, 12'hB88, 12'hD99, 12'hC88, 12'hB87, 12'hB88, 12'hA77, 12'hB88, 12'hB98, 12'hB87, 12'hB77, 12'hC88, 12'hC88, 12'hB77, 12'hB87, 12'hB77, 12'hA77, 12'hA76, 12'hA66, 12'hA66, 12'h865, 12'h855, 12'h855, 12'h754, 12'h744, 12'h644, 12'h644, 12'h644, 12'h543, 12'h644, 12'h644, 12'h644, 12'h543, 12'h533, 12'h433, 12'h332, 12'h543, 12'h433, 12'h433, 12'h333, 12'h332, 12'h322, 12'h222, 12'h221, 12'h221, 12'h221, 12'h211, 12'h111, 12'h221, 12'h222, 12'h666, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCB, 12'hBBC, 12'hCBB, 12'hCCB, 12'hBBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hCCC, 12'hBCB, 12'hCBB, 12'hCCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCDC, 12'hCCC, 12'hBBB, 12'hBAB, 12'h999, 12'h778, 12'h667, 12'h999, 12'h889, 12'h878, 12'h777, 12'h989, 12'h989, 12'h99A, 12'h777, 12'h878, 12'h878, 12'h878, 12'h888, 12'h656, 12'h655, 12'h322, 12'h644, 12'hB88, 12'hD98, 12'hD98, 12'hB77, 12'hC87, 12'hD88, 12'hD98, 12'hB77, 12'h966, 12'h976, 12'hA77, 12'h966, 12'h866, 12'h866, 12'h865, 12'h755, 12'h745, 12'h644, 12'h644, 12'h644, 12'h655, 12'h755, 12'h644, 12'h655, 12'h654, 12'h644, 12'h654, 12'h644, 12'h755, 12'h755, 12'h866, 12'h976, 12'h866, 12'h966, 12'h977, 12'hB88, 12'hC99, 12'hC88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hA77, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hA77, 12'hC88, 12'hB77, 12'hA66, 12'hA76, 12'hA66, 12'hA66, 12'h965, 12'h965, 12'h855, 12'h854, 12'h754, 12'h644, 12'h644, 12'h643, 12'h644, 12'h543, 12'h533, 12'h544, 12'h543, 12'h533, 12'h543, 12'h433, 12'h443, 12'h333, 12'h544, 12'h333, 12'h332, 12'h333, 12'h322, 12'h222, 12'h222, 12'h221, 12'h221, 12'h111, 12'h111, 12'h221, 12'h222, 12'h222, 12'hCBC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCB, 12'hCBC, 12'hBCB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hCBC, 12'hCCB, 12'hBBB, 12'hCCC, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCC, 12'hCCC, 12'hCBB, 12'hBCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBBB, 12'hAAA, 12'h777, 12'h878, 12'h767, 12'h99A, 12'h999, 12'h888, 12'h999, 12'h989, 12'h889, 12'h878, 12'h878, 12'h777, 12'h878, 12'h777, 12'h888, 12'h878, 12'h767, 12'h544, 12'h322, 12'h876, 12'hB88, 12'hDA8, 12'hC98, 12'hB87, 12'hC87, 12'hD98, 12'hD87, 12'hB77, 12'h966, 12'h976, 12'h976, 12'h866, 12'h967, 12'h866, 12'h755, 12'h755, 12'h755, 12'h755, 12'h755, 12'h755, 12'h644, 12'h644, 12'h755, 12'h644, 12'h544, 12'h544, 12'h544, 12'h644, 12'h654, 12'h865, 12'h966, 12'h977, 12'hA88, 12'hA87, 12'hB88, 12'hA78, 12'hB98, 12'hC88, 12'hC88, 12'hB88, 12'hB88, 12'hB88, 12'hA77, 12'hB88, 12'hB88, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hB77, 12'hA76, 12'hA77, 12'hA77, 12'hA66, 12'h966, 12'h854, 12'h855, 12'h855, 12'h754, 12'h755, 12'h744, 12'h644, 12'h533, 12'h544, 12'h544, 12'h533, 12'h543, 12'h544, 12'h433, 12'h433, 12'h443, 12'h433, 12'h544, 12'h443, 12'h433, 12'h433, 12'h232, 12'h222, 12'h222, 12'h221, 12'h211, 12'h111, 12'h111, 12'h121, 12'h222, 12'h222, 12'h777, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDCC, 12'hCCD, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hBCB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBCB, 12'hCCC, 12'hCCC, 12'hBCB, 12'hBCC, 12'hBBB, 12'hAAA, 12'hAAA, 12'h99A, 12'h999, 12'hAAA, 12'hAAB, 12'h989, 12'h777, 12'h444, 12'h777, 12'h888, 12'h989, 12'h889, 12'h878, 12'hAAA, 12'h888, 12'h878, 12'h777, 12'h777, 12'h778, 12'h889, 12'h778, 12'h777, 12'h766, 12'h333, 12'h432, 12'h976, 12'hB87, 12'hD98, 12'hC87, 12'hB76, 12'hC87, 12'hD87, 12'hC87, 12'hB77, 12'h966, 12'h866, 12'h866, 12'h866, 12'h866, 12'h866, 12'h866, 12'h755, 12'h755, 12'h754, 12'h754, 12'h755, 12'h655, 12'h654, 12'h655, 12'h644, 12'h755, 12'h544, 12'h655, 12'h644, 12'h655, 12'h766, 12'h866, 12'h966, 12'hA88, 12'h977, 12'hB88, 12'hA87, 12'hC99, 12'hC98, 12'hB88, 12'hB87, 12'hA87, 12'hB87, 12'hA77, 12'hA77, 12'hA77, 12'h966, 12'h966, 12'hB77, 12'hA76, 12'hA77, 12'hA76, 12'hA77, 12'h966, 12'h855, 12'h865, 12'h865, 12'h755, 12'h754, 12'h855, 12'h744, 12'h544, 12'h544, 12'h544, 12'h544, 12'h543, 12'h433, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h322, 12'h222, 12'h222, 12'h221, 12'h121, 12'h111, 12'h111, 12'h222, 12'h222, 12'h333, 12'h889, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDED, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDD, 12'hDDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCCC, 12'hCCB, 12'hCBC, 12'hCBB, 12'hBCB, 12'hCBC, 12'hBBB, 12'hBCB, 12'hCBC, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'hBBB, 12'hBBB, 12'hA9A, 12'h888, 12'h889, 12'h989, 12'h989, 12'h888, 12'h878, 12'h889, 12'hBBB, 12'hBAB, 12'h999, 12'h555, 12'h444, 12'h656, 12'h888, 12'h667, 12'h767, 12'h888, 12'h878, 12'h888, 12'h666, 12'h778, 12'h767, 12'h666, 12'h777, 12'h767, 12'h878, 12'h767, 12'h655, 12'h333, 12'h533, 12'h976, 12'hC87, 12'hC98, 12'hC87, 12'hB77, 12'hC87, 12'hD98, 12'hC87, 12'hB87, 12'hA77, 12'h866, 12'h866, 12'h866, 12'h866, 12'h766, 12'h755, 12'h655, 12'h644, 12'h655, 12'h755, 12'h755, 12'h755, 12'h755, 12'h645, 12'h544, 12'h644, 12'h544, 12'h544, 12'h544, 12'h655, 12'h766, 12'h755, 12'h866, 12'h977, 12'hA76, 12'hB87, 12'hA77, 12'hB77, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'h865, 12'h966, 12'h977, 12'h966, 12'h966, 12'hA77, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h966, 12'h966, 12'h866, 12'h866, 12'h744, 12'h744, 12'h855, 12'h755, 12'h533, 12'h543, 12'h543, 12'h533, 12'h534, 12'h433, 12'h433, 12'h332, 12'h332, 12'h433, 12'h333, 12'h332, 12'h322, 12'h232, 12'h222, 12'h221, 12'h221, 12'h111, 12'h111, 12'h221, 12'h221, 12'h222, 12'h666, 12'hCCD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hEDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDCD, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBB, 12'hCBC, 12'hCCB, 12'hCBB, 12'hCBC, 12'hBCB, 12'hCBB, 12'hBBC, 12'hCCB, 12'hCBB, 12'hCBC, 12'hBCB, 12'hCBB, 12'hBCC, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB,
		12'h989, 12'h888, 12'h989, 12'h888, 12'h878, 12'h777, 12'h878, 12'h666, 12'h555, 12'h445, 12'h99A, 12'hA9A, 12'hAAA, 12'h989, 12'h666, 12'h444, 12'h555, 12'h545, 12'h445, 12'h556, 12'h556, 12'h889, 12'h656, 12'h777, 12'h889, 12'h767, 12'h767, 12'h878, 12'h777, 12'h767, 12'h555, 12'h544, 12'h433, 12'h544, 12'h966, 12'hB87, 12'hC87, 12'hB77, 12'hB76, 12'hC87, 12'hD98, 12'hD87, 12'hC87, 12'hA76, 12'h866, 12'h866, 12'h866, 12'h766, 12'h866, 12'h755, 12'h645, 12'h655, 12'h644, 12'h754, 12'h755, 12'h755, 12'h754, 12'h644, 12'h644, 12'h655, 12'h655, 12'h544, 12'h644, 12'h655, 12'h655, 12'h866, 12'hA78, 12'h966, 12'hA87, 12'hA76, 12'hB87, 12'hB77, 12'h976, 12'h865, 12'h966, 12'hA76, 12'h976, 12'h855, 12'h866, 12'h855, 12'h876, 12'h866, 12'h865, 12'h865, 12'h866, 12'h855, 12'h755, 12'h855, 12'h755, 12'h644, 12'h654, 12'h644, 12'h544, 12'h433, 12'h544, 12'h544, 12'h433, 12'h443, 12'h333, 12'h333, 12'h322, 12'h332, 12'h333, 12'h322, 12'h333, 12'h222, 12'h222, 12'h221, 12'h111, 12'h221, 12'h111, 12'h221, 12'h222, 12'h222, 12'h888, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCCD, 12'hDDC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hBCC, 12'hBCB, 12'hBBB, 12'hBCC, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hBBB,
		12'h888, 12'h767, 12'h767, 12'h667, 12'h444, 12'h444, 12'h555, 12'h334, 12'h333, 12'h555, 12'h99A, 12'hAAA, 12'h989, 12'h889, 12'h555, 12'h333, 12'h334, 12'h444, 12'h444, 12'h556, 12'h767, 12'h666, 12'h778, 12'h667, 12'h667, 12'h777, 12'h767, 12'h888, 12'h667, 12'h777, 12'h556, 12'h545, 12'h433, 12'h432, 12'h644, 12'h966, 12'hA76, 12'hB87, 12'hB77, 12'hB76, 12'hC87, 12'hC88, 12'hC87, 12'hB87, 12'hB77, 12'h866, 12'h766, 12'h756, 12'h866, 12'h766, 12'h766, 12'h655, 12'h645, 12'h755, 12'h755, 12'h855, 12'h655, 12'h755, 12'h755, 12'h655, 12'h644, 12'h644, 12'h544, 12'h655, 12'h544, 12'h644, 12'h877, 12'h765, 12'h866, 12'h866, 12'h966, 12'hA76, 12'h866, 12'h966, 12'h866, 12'h855, 12'h755, 12'h755, 12'h754, 12'h866, 12'h755, 12'h866, 12'h855, 12'h865, 12'h744, 12'h644, 12'h644, 12'h755, 12'h543, 12'h543, 12'h544, 12'h534, 12'h433, 12'h544, 12'h433, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h333, 12'h222, 12'h222, 12'h221, 12'h222, 12'h221, 12'h111, 12'h121, 12'h212, 12'h111, 12'h222, 12'h222, 12'h333, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDED, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCCC, 12'hCCD, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCCC, 12'hCBB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCBC, 12'hBCB, 12'hCBB, 12'hBBC, 12'hBCB, 12'hCBB, 12'hBBC, 12'hBBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBBB,
		12'h556, 12'h555, 12'h666, 12'h656, 12'h334, 12'h333, 12'h334, 12'h556, 12'h778, 12'h767, 12'h767, 12'hAAA, 12'h99A, 12'h99A, 12'h989, 12'h777, 12'h333, 12'h333, 12'h333, 12'h444, 12'h667, 12'h667, 12'h778, 12'h666, 12'h556, 12'h767, 12'h445, 12'h778, 12'h667, 12'h656, 12'h767, 12'h444, 12'h445, 12'h433, 12'h432, 12'h543, 12'h855, 12'hA76, 12'hB87, 12'hB77, 12'hA76, 12'hB87, 12'hC88, 12'hB87, 12'hA77, 12'hB77, 12'h977, 12'h855, 12'h755, 12'h766, 12'h755, 12'h755, 12'h655, 12'h544, 12'h644, 12'h655, 12'h644, 12'h755, 12'h644, 12'h755, 12'h755, 12'h644, 12'h644, 12'h544, 12'h655, 12'h544, 12'h544, 12'h644, 12'h766, 12'h755, 12'h865, 12'h866, 12'h966, 12'h866, 12'h654, 12'h644, 12'h755, 12'h754, 12'h755, 12'h644, 12'h644, 12'h755, 12'h644, 12'h755, 12'h533, 12'h644, 12'h654, 12'h543, 12'h543, 12'h433, 12'h433, 12'h322, 12'h332, 12'h332, 12'h321, 12'h322, 12'h222, 12'h322, 12'h222, 12'h221, 12'h322, 12'h222, 12'h222, 12'h211, 12'h111, 12'h121, 12'h211, 12'h111, 12'h221, 12'h221, 12'h222, 12'h222, 12'h222, 12'h899, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCCB, 12'hBBB, 12'hCCC, 12'hCCB, 12'hBBC, 12'hCBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hCCB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hCBB, 12'hBCB, 12'hBBB, 12'hBCB, 12'hCCB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hCBB,
		12'h667, 12'h666, 12'h556, 12'h555, 12'h445, 12'h556, 12'h888, 12'h878, 12'h767, 12'h667, 12'h666, 12'h889, 12'hBAB, 12'h999, 12'h989, 12'h989, 12'h556, 12'h323, 12'h333, 12'h334, 12'h334, 12'h444, 12'h656, 12'h656, 12'h556, 12'h767, 12'h667, 12'h555, 12'h777, 12'h767, 12'h555, 12'h445, 12'h666, 12'h333, 12'h333, 12'h432, 12'h533, 12'h855, 12'hA76, 12'hB87, 12'hB77, 12'hA66, 12'hB77, 12'hD98, 12'hD88, 12'hB87, 12'hB87, 12'hB88, 12'h856, 12'h755, 12'h755, 12'h855, 12'h765, 12'h655, 12'h644, 12'h544, 12'h644, 12'h754, 12'h754, 12'h644, 12'h755, 12'h644, 12'h654, 12'h644, 12'h655, 12'h544, 12'h544, 12'h544, 12'h544, 12'h655, 12'h655, 12'h655, 12'h755, 12'h654, 12'h644, 12'h644, 12'h433, 12'h543, 12'h655, 12'h543, 12'h544, 12'h433, 12'h544, 12'h544, 12'h543, 12'h543, 12'h422, 12'h433, 12'h322, 12'h433, 12'h222, 12'h333, 12'h322, 12'h433, 12'h222, 12'h221, 12'h211, 12'h211, 12'h121, 12'h222, 12'h222, 12'h221, 12'h111, 12'h111, 12'h221, 12'h111, 12'h111, 12'h121, 12'h211, 12'h111, 12'h222, 12'h222, 12'h333, 12'hDCD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hCDC, 12'hCCD, 12'hDCD, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBCC, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBBC, 12'hCBB, 12'hCBC, 12'hBBC, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hCBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBCB, 12'hCBC, 12'hCCB, 12'hCCC,
		12'h555, 12'h545, 12'h445, 12'h667, 12'h778, 12'h999, 12'h878, 12'h767, 12'h666, 12'h555, 12'h677, 12'h778, 12'h99A, 12'hAAA, 12'hAAA, 12'hA9A, 12'h989, 12'h777, 12'h444, 12'h333, 12'h333, 12'h334, 12'h555, 12'h556, 12'h555, 12'h556, 12'h656, 12'h767, 12'h667, 12'h777, 12'h666, 12'h555, 12'h656, 12'h545, 12'h434, 12'h433, 12'h432, 12'h533, 12'h855, 12'hA76, 12'hC87, 12'hC87, 12'hA66, 12'hB77, 12'hD87, 12'hC87, 12'hC87, 12'hB87, 12'hB87, 12'h967, 12'h655, 12'h755, 12'h755, 12'h655, 12'h655, 12'h655, 12'h544, 12'h644, 12'h644, 12'h655, 12'h644, 12'h655, 12'h755, 12'h644, 12'h544, 12'h644, 12'h544, 12'h645, 12'h645, 12'h534, 12'h433, 12'h434, 12'h544, 12'h544, 12'h444, 12'h433, 12'h433, 12'h323, 12'h333, 12'h333, 12'h322, 12'h333, 12'h333, 12'h433, 12'h444, 12'h322, 12'h322, 12'h212, 12'h222, 12'h221, 12'h222, 12'h222, 12'h211, 12'h111, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h110, 12'h111, 12'h111, 12'h221, 12'h111, 12'h111, 12'h221, 12'h121, 12'h222, 12'h111, 12'h221, 12'h666, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hCDD, 12'hDCC, 12'hCCC, 12'hCDD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCCC, 12'hCBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBBB, 12'hCCB, 12'hBCB, 12'hCBC, 12'hCBB, 12'hBCB, 12'hCBB, 12'hBBC, 12'hBCB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBCC, 12'hCCB, 12'hCCB,
		12'h667, 12'h667, 12'h777, 12'h777, 12'h878, 12'h555, 12'h556, 12'h667, 12'h667, 12'h878, 12'h889, 12'h767, 12'h778, 12'h989, 12'hAAB, 12'hAAB, 12'h888, 12'hAAA, 12'h989, 12'h888, 12'h667, 12'h656, 12'h666, 12'h556, 12'h667, 12'h767, 12'h667, 12'h667, 12'h667, 12'h667, 12'h556, 12'h656, 12'h656, 12'h444, 12'h445, 12'h434, 12'h433, 12'h432, 12'h543, 12'h955, 12'hA66, 12'hB76, 12'hC87, 12'hA76, 12'hA76, 12'hB77, 12'hB77, 12'hA77, 12'hB87, 12'hB87, 12'h976, 12'h866, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h543, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h654, 12'h644, 12'h544, 12'h544, 12'h544, 12'h433, 12'h333, 12'h322, 12'h222, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h221, 12'h212, 12'h211, 12'h121, 12'h222, 12'h111, 12'h111, 12'h211, 12'h111, 12'h211, 12'h111, 12'h111, 12'h111, 12'h110, 12'h111, 12'h110, 12'h110, 12'h110, 12'h110, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h221, 12'h211, 12'h111, 12'h211, 12'h221, 12'h222, 12'hAAB, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hCCD, 12'hDDC, 12'hCDD, 12'hDCC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBBC, 12'hCCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCBB, 12'hBBB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBBB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCCC, 12'hBBB, 12'hBCB, 12'hCCC, 12'hBBB, 12'hBBB, 12'hCCB, 12'hBBB, 12'hBCB, 12'hCCB, 12'hBBC, 12'hCCB, 12'hCCB, 12'hCBB,
		12'h767, 12'h888, 12'h666, 12'h656, 12'h666, 12'h888, 12'h989, 12'h767, 12'h666, 12'h444, 12'h333, 12'h222, 12'h334, 12'h778, 12'h878, 12'h889, 12'h889, 12'h99A, 12'h989, 12'hA9A, 12'h889, 12'hAAA, 12'hAAA, 12'hAAA, 12'hCBC, 12'hA99, 12'h555, 12'h555, 12'h666, 12'h656, 12'h555, 12'h556, 12'h555, 12'h556, 12'h556, 12'h445, 12'h445, 12'h433, 12'h432, 12'h644, 12'h855, 12'hA65, 12'hC87, 12'hC87, 12'hB87, 12'h965, 12'h966, 12'hA77, 12'hB77, 12'hB77, 12'hB77, 12'hA77, 12'h966, 12'h655, 12'h544, 12'h433, 12'h544, 12'h644, 12'h544, 12'h543, 12'h543, 12'h544, 12'h544, 12'h543, 12'h644, 12'h544, 12'h644, 12'h655, 12'h644, 12'h544, 12'h544, 12'h544, 12'h544, 12'h433, 12'h433, 12'h322, 12'h332, 12'h322, 12'h221, 12'h211, 12'h211, 12'h211, 12'h211, 12'h221, 12'h111, 12'h110, 12'h111, 12'h111, 12'h111, 12'h211, 12'h111, 12'h110, 12'h111, 12'h110, 12'h110, 12'h110, 12'h111, 12'h111, 12'h110, 12'h111, 12'h110, 12'h110, 12'h111, 12'h110, 12'h110, 12'h111, 12'h211, 12'h121, 12'h111, 12'h222, 12'h222, 12'h333, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDDD, 12'hCCC, 12'hDCD, 12'hCDC, 12'hCCC, 12'hDCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hBCC, 12'hCCB, 12'hBBB, 12'hBCC, 12'hCCB, 12'hBBB, 12'hCCC, 12'hBCB, 12'hBBB, 12'hCBC, 12'hBCB, 12'hCBC, 12'hCCC, 12'hCBB, 12'hBBC, 12'hCCB, 12'hBBB, 12'hBBC, 12'hCCB, 12'hBCB, 12'hCBC, 12'hCCB, 12'hBBB, 12'hCBC, 12'hBCB, 12'hBCC, 12'hCBB, 12'hCCB, 12'hCCB,
		12'h656, 12'h777, 12'h888, 12'h778, 12'h767, 12'h445, 12'h334, 12'h223, 12'h333, 12'h333, 12'h333, 12'h555, 12'h334, 12'h444, 12'h667, 12'h666, 12'h767, 12'h556, 12'h667, 12'h667, 12'h667, 12'h889, 12'h99A, 12'hBBB, 12'h777, 12'h555, 12'h555, 12'h555, 12'h656, 12'h555, 12'h444, 12'h667, 12'h556, 12'h656, 12'h545, 12'h555, 12'h545, 12'h434, 12'h322, 12'h432, 12'h644, 12'h855, 12'hB76, 12'hC87, 12'hC87, 12'hC87, 12'hA76, 12'h965, 12'h866, 12'hB77, 12'hB77, 12'hB77, 12'h976, 12'h866, 12'h866, 12'h766, 12'h544, 12'h433, 12'h433, 12'h533, 12'h544, 12'h433, 12'h433, 12'h433, 12'h544, 12'h544, 12'h644, 12'h644, 12'h644, 12'h644, 12'h433, 12'h533, 12'h543, 12'h433, 12'h534, 12'h433, 12'h433, 12'h433, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h211, 12'h211, 12'h211, 12'h211, 12'h110, 12'h110, 12'h111, 12'h111, 12'h110, 12'h110, 12'h110, 12'h100, 12'h110, 12'h100, 12'h010, 12'h110, 12'h111, 12'h110, 12'h111, 12'h110, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h221, 12'h222, 12'h222, 12'h999, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDD, 12'hDDC, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCBC, 12'hCBC, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hCCB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBCB, 12'hBCC, 12'hBCC, 12'hBCC, 12'hCBC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC,
		12'h555, 12'h666, 12'h445, 12'h444, 12'h333, 12'h333, 12'h434, 12'h444, 12'h334, 12'h333, 12'h334, 12'h444, 12'h334, 12'h444, 12'h556, 12'h777, 12'h656, 12'h656, 12'h556, 12'h778, 12'h878, 12'h888, 12'h767, 12'h767, 12'h555, 12'h444, 12'h333, 12'h444, 12'h444, 12'h555, 12'h444, 12'h445, 12'h445, 12'h555, 12'h444, 12'h445, 12'h444, 12'h444, 12'h333, 12'h213, 12'h323, 12'h543, 12'h855, 12'hA76, 12'hB76, 12'hC87, 12'hC87, 12'hB77, 12'h966, 12'h865, 12'h966, 12'hA66, 12'h966, 12'hA76, 12'h966, 12'h966, 12'h866, 12'h755, 12'h644, 12'h544, 12'h433, 12'h433, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h221, 12'h211, 12'h211, 12'h211, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h110, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h221, 12'h221, 12'h222, 12'h222, 12'h222, 12'h555, 12'h999, 12'hCDC, 12'hDDD, 12'hDDD, 12'hDDD, 12'hCDC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCBB, 12'hCBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBBB, 12'hBCB, 12'hBCB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCB, 12'hCCB, 12'hCCC, 12'hCCC, 12'hBCC, 12'hBCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC,};

	assign rgb_colour = array[160*v_count_n+h_count_n];
endmodule