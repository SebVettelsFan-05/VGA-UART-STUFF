module image_rom (
	input logic [9:0] v_count,
	input logic [9:0] h_count,
	output logic [11:0] rgb_colour
);
	logic [9:0] v_count_n;
	logic [9:0] h_count_n;
	assign v_count_n = v_count >> 2;
	assign h_count_n = h_count >> 2;

	logic [11:0] array[0:19199] = '{
		12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h455, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444,
		12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h455, 12'h445, 12'h445, 12'h455, 12'h445, 12'h554, 12'h455, 12'h445, 12'h554, 12'h455, 12'h545, 12'h455, 12'h445, 12'h444, 12'h445, 12'h455, 12'h544, 12'h555, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444,
		12'h444, 12'h445, 12'h434, 12'h444, 12'h444, 12'h434, 12'h445, 12'h444, 12'h434, 12'h444, 12'h444, 12'h435, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h555, 12'h554, 12'h445, 12'h554, 12'h545, 12'h444, 12'h455, 12'h545, 12'h544, 12'h455, 12'h554, 12'h445, 12'h555, 12'h454, 12'h444, 12'h555, 12'h444, 12'h454, 12'h555, 12'h555, 12'h444, 12'h555, 12'h454, 12'h445, 12'h454, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444,
		12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h435, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h554, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h454, 12'h544, 12'h455, 12'h544, 12'h445, 12'h454, 12'h554, 12'h445, 12'h454, 12'h544, 12'h455, 12'h445, 12'h544, 12'h455, 12'h444, 12'h545, 12'h444, 12'h444, 12'h545, 12'h445, 12'h444, 12'h555, 12'h445, 12'h444, 12'h554, 12'h545, 12'h444, 12'h554, 12'h445, 12'h444, 12'h554, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444,
		12'h444, 12'h445, 12'h444, 12'h444, 12'h435, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h544, 12'h555, 12'h444, 12'h445, 12'h455, 12'h445, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h455, 12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h554, 12'h445, 12'h454, 12'h545, 12'h455, 12'h554, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h444, 12'h455, 12'h545, 12'h455, 12'h455, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h544, 12'h455, 12'h554, 12'h444, 12'h445, 12'h444,
		12'h444, 12'h445, 12'h444, 12'h444, 12'h434, 12'h444, 12'h445, 12'h434, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h545, 12'h444, 12'h444, 12'h545, 12'h445, 12'h444, 12'h544, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h445, 12'h444, 12'h555, 12'h445, 12'h444, 12'h445, 12'h444, 12'h454, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h455, 12'h445, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h455, 12'h455, 12'h444, 12'h455, 12'h454, 12'h445, 12'h454, 12'h444, 12'h445, 12'h455, 12'h544, 12'h445, 12'h455, 12'h554, 12'h555, 12'h444, 12'h554, 12'h555, 12'h444, 12'h444, 12'h555, 12'h445, 12'h554, 12'h455, 12'h545, 12'h445, 12'h455, 12'h545, 12'h444, 12'h454, 12'h555, 12'h445, 12'h554, 12'h554, 12'h445, 12'h554, 12'h455, 12'h445, 12'h555, 12'h455, 12'h444, 12'h445, 12'h455, 12'h544, 12'h445, 12'h445, 12'h444, 12'h444,
		12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h544, 12'h445, 12'h445, 12'h544, 12'h445, 12'h445, 12'h444, 12'h545, 12'h445, 12'h454, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h444, 12'h445, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h455, 12'h545, 12'h455, 12'h545, 12'h555, 12'h455, 12'h444, 12'h545, 12'h455, 12'h445, 12'h455, 12'h454, 12'h445, 12'h455, 12'h455, 12'h444, 12'h445, 12'h455, 12'h444, 12'h545, 12'h455, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h455, 12'h545, 12'h554, 12'h555, 12'h545, 12'h555, 12'h554, 12'h445, 12'h555, 12'h445, 12'h554, 12'h445, 12'h444, 12'h555, 12'h444, 12'h445, 12'h555, 12'h445, 12'h445, 12'h554, 12'h455, 12'h545, 12'h454, 12'h445, 12'h555, 12'h444, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h445, 12'h555, 12'h545, 12'h455, 12'h545, 12'h455, 12'h545, 12'h554, 12'h455, 12'h545, 12'h554, 12'h555, 12'h445, 12'h554, 12'h545, 12'h444, 12'h454, 12'h545, 12'h444, 12'h445,
		12'h444, 12'h444, 12'h444, 12'h445, 12'h434, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h454, 12'h544, 12'h445, 12'h454, 12'h445, 12'h544, 12'h454, 12'h445, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h455, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h455, 12'h445, 12'h444, 12'h555, 12'h555, 12'h444, 12'h445, 12'h555, 12'h555, 12'h444, 12'h445, 12'h545, 12'h444, 12'h545, 12'h445, 12'h555, 12'h555, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h454, 12'h555, 12'h545, 12'h445, 12'h455, 12'h555, 12'h445, 12'h444, 12'h555, 12'h545, 12'h444, 12'h555, 12'h445, 12'h454, 12'h544, 12'h455, 12'h454, 12'h544, 12'h445, 12'h454, 12'h545, 12'h445, 12'h455, 12'h545, 12'h554, 12'h455, 12'h545, 12'h444, 12'h555, 12'h455, 12'h554, 12'h555, 12'h455, 12'h554, 12'h545, 12'h454, 12'h555, 12'h455, 12'h545, 12'h455, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h545, 12'h555, 12'h455, 12'h445, 12'h554, 12'h444, 12'h455, 12'h555,
		12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h455, 12'h454, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h454, 12'h444, 12'h444, 12'h455, 12'h555, 12'h544, 12'h444, 12'h444, 12'h544, 12'h444, 12'h555, 12'h444, 12'h444, 12'h544, 12'h555, 12'h444, 12'h544, 12'h554, 12'h444, 12'h444, 12'h444, 12'h544, 12'h444, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h433, 12'h444, 12'h544, 12'h444, 12'h433, 12'h444, 12'h434, 12'h444, 12'h434, 12'h444, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h444, 12'h333, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h554, 12'h555, 12'h455, 12'h455, 12'h544, 12'h455, 12'h555, 12'h445, 12'h455, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h455, 12'h544, 12'h444, 12'h555, 12'h544, 12'h545, 12'h455, 12'h545, 12'h545, 12'h545,
		12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h545, 12'h445, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h544, 12'h444, 12'h544, 12'h455, 12'h444, 12'h545, 12'h455, 12'h444, 12'h545, 12'h455, 12'h445, 12'h554, 12'h445, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h454, 12'h445, 12'h444, 12'h445, 12'h445, 12'h544, 12'h444, 12'h444, 12'h444, 12'h555, 12'h554, 12'h444, 12'h444, 12'h545, 12'h544, 12'h554, 12'h555, 12'h555, 12'h555, 12'h544, 12'h444, 12'h555, 12'h555, 12'h544, 12'h544, 12'h555, 12'h655, 12'h656, 12'h555, 12'h555, 12'h555, 12'h555, 12'h544, 12'h555, 12'h655, 12'h655, 12'h666, 12'h544, 12'h544, 12'h544, 12'h444, 12'h434, 12'h444, 12'h544, 12'h434, 12'h434, 12'h433, 12'h444, 12'h444, 12'h444, 12'h333, 12'h333, 12'h433, 12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h444, 12'h544, 12'h455, 12'h544, 12'h445, 12'h455, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h455, 12'h554, 12'h555, 12'h555, 12'h555, 12'h445, 12'h455, 12'h554, 12'h444, 12'h555, 12'h545, 12'h444, 12'h445,
		12'h444, 12'h445, 12'h444, 12'h445, 12'h545, 12'h444, 12'h545, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h455, 12'h444, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h544, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h445, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h545, 12'h454, 12'h544, 12'h544, 12'h444, 12'h544, 12'h555, 12'h555, 12'h545, 12'h444, 12'h555, 12'h544, 12'h444, 12'h545, 12'h555, 12'h544, 12'h545, 12'h655, 12'h555, 12'h545, 12'h544, 12'h544, 12'h444, 12'h444, 12'h444, 12'h545, 12'h545, 12'h555, 12'h555, 12'h545, 12'h655, 12'h656, 12'h555, 12'h655, 12'h555, 12'h555, 12'h555, 12'h545, 12'h444, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h433, 12'h333, 12'h333, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h444, 12'h445, 12'h555, 12'h454, 12'h555, 12'h555, 12'h454, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h445, 12'h554, 12'h455, 12'h444, 12'h544,
		12'h445, 12'h444, 12'h545, 12'h444, 12'h445, 12'h545, 12'h444, 12'h445, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h544, 12'h444, 12'h444, 12'h544, 12'h445, 12'h544, 12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h554, 12'h445, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h454, 12'h445, 12'h444, 12'h454, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h445, 12'h454, 12'h445, 12'h445, 12'h454, 12'h444, 12'h445, 12'h544, 12'h444, 12'h454, 12'h444, 12'h555, 12'h555, 12'h655, 12'h656, 12'h655, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h655, 12'h655, 12'h666, 12'h666, 12'h655, 12'h545, 12'h555, 12'h555, 12'h555, 12'h655, 12'h655, 12'h655, 12'h555, 12'h544, 12'h544, 12'h544, 12'h444, 12'h544, 12'h444, 12'h444, 12'h555, 12'h655, 12'h656, 12'h555, 12'h544, 12'h544, 12'h544, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h544, 12'h434, 12'h333, 12'h333, 12'h333, 12'h223, 12'h333, 12'h444, 12'h445, 12'h545, 12'h555, 12'h555, 12'h445, 12'h555, 12'h545, 12'h455, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h545, 12'h545, 12'h455, 12'h544, 12'h545, 12'h545,
		12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h545, 12'h444, 12'h445, 12'h545, 12'h444, 12'h445, 12'h444, 12'h454, 12'h545, 12'h454, 12'h445, 12'h544, 12'h455, 12'h445, 12'h544, 12'h455, 12'h444, 12'h444, 12'h445, 12'h445, 12'h544, 12'h455, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h455, 12'h445, 12'h444, 12'h455, 12'h444, 12'h444, 12'h444, 12'h455, 12'h555, 12'h444, 12'h555, 12'h544, 12'h444, 12'h655, 12'h666, 12'h767, 12'h777, 12'h777, 12'h766, 12'h666, 12'h655, 12'h555, 12'h544, 12'h443, 12'h444, 12'h444, 12'h544, 12'h555, 12'h555, 12'h554, 12'h555, 12'h544, 12'h544, 12'h443, 12'h433, 12'h433, 12'h434, 12'h544, 12'h554, 12'h655, 12'h666, 12'h666, 12'h655, 12'h555, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h555, 12'h554, 12'h554, 12'h544, 12'h544, 12'h545, 12'h544, 12'h444, 12'h433, 12'h433, 12'h333, 12'h433, 12'h444, 12'h555, 12'h444, 12'h433, 12'h333, 12'h333, 12'h333, 12'h323, 12'h222, 12'h333, 12'h333, 12'h444, 12'h555, 12'h554, 12'h445, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h545, 12'h455, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h554, 12'h545, 12'h555, 12'h545, 12'h545,
		12'h444, 12'h445, 12'h444, 12'h445, 12'h545, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h544, 12'h444, 12'h444, 12'h445, 12'h444, 12'h554, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h445, 12'h454, 12'h444, 12'h444, 12'h544, 12'h444, 12'h444, 12'h545, 12'h444, 12'h445, 12'h555, 12'h455, 12'h444, 12'h444, 12'h444, 12'h444, 12'h555, 12'h666, 12'h877, 12'h888, 12'h777, 12'h776, 12'h776, 12'h766, 12'h666, 12'h666, 12'h766, 12'h766, 12'h655, 12'h554, 12'h555, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h555, 12'h544, 12'h544, 12'h544, 12'h545, 12'h544, 12'h544, 12'h655, 12'h655, 12'h655, 12'h666, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h655, 12'h655, 12'h555, 12'h654, 12'h544, 12'h545, 12'h544, 12'h544, 12'h444, 12'h444, 12'h544, 12'h545, 12'h545, 12'h444, 12'h544, 12'h444, 12'h333, 12'h333, 12'h444, 12'h333, 12'h333, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h323, 12'h222, 12'h333, 12'h444, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h455, 12'h445, 12'h545, 12'h555, 12'h455, 12'h445, 12'h555, 12'h555, 12'h445, 12'h545,
		12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h545, 12'h455, 12'h444, 12'h545, 12'h445, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h454, 12'h444, 12'h445, 12'h444, 12'h455, 12'h444, 12'h444, 12'h454, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h555, 12'h666, 12'h877, 12'h888, 12'h877, 12'h888, 12'h888, 12'h777, 12'h665, 12'h655, 12'h766, 12'h877, 12'h776, 12'h665, 12'h655, 12'h666, 12'h655, 12'h665, 12'h656, 12'h655, 12'h554, 12'h655, 12'h655, 12'h544, 12'h544, 12'h655, 12'h655, 12'h544, 12'h544, 12'h555, 12'h555, 12'h544, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h766, 12'h766, 12'h766, 12'h655, 12'h544, 12'h544, 12'h544, 12'h544, 12'h434, 12'h433, 12'h333, 12'h333, 12'h434, 12'h434, 12'h444, 12'h444, 12'h545, 12'h444, 12'h222, 12'h433, 12'h333, 12'h323, 12'h333, 12'h434, 12'h333, 12'h322, 12'h222, 12'h223, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h544, 12'h555, 12'h545, 12'h444, 12'h555, 12'h555,
		12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h544, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h445, 12'h444, 12'h544, 12'h445, 12'h444, 12'h545, 12'h455, 12'h545, 12'h444, 12'h444, 12'h555, 12'h444, 12'h544, 12'h545, 12'h555, 12'h777, 12'h988, 12'h888, 12'h878, 12'h777, 12'h776, 12'h766, 12'h766, 12'h766, 12'h777, 12'h877, 12'h777, 12'h766, 12'h766, 12'h766, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h766, 12'h766, 12'h766, 12'h876, 12'h877, 12'h766, 12'h766, 12'h766, 12'h766, 12'h766, 12'h765, 12'h766, 12'h766, 12'h755, 12'h655, 12'h654, 12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h554, 12'h544, 12'h434, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h322, 12'h323, 12'h444, 12'h433, 12'h434, 12'h333, 12'h333, 12'h333, 12'h323, 12'h333, 12'h323, 12'h332, 12'h322, 12'h222, 12'h222, 12'h323, 12'h333, 12'h444, 12'h445, 12'h545, 12'h445, 12'h455, 12'h556, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h554, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555,
		12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h444, 12'h454, 12'h544, 12'h545, 12'h444, 12'h444, 12'h555, 12'h544, 12'h666, 12'h777, 12'h777, 12'h666, 12'h767, 12'h656, 12'h777, 12'h777, 12'h666, 12'h655, 12'h766, 12'h766, 12'h666, 12'h655, 12'h655, 12'h766, 12'h655, 12'h654, 12'h655, 12'h766, 12'h766, 12'h765, 12'h655, 12'h655, 12'h755, 12'h755, 12'h755, 12'h766, 12'h755, 12'h756, 12'h766, 12'h866, 12'h866, 12'h877, 12'h988, 12'h877, 12'h866, 12'h877, 12'h876, 12'h866, 12'h766, 12'h765, 12'h755, 12'h755, 12'h655, 12'h654, 12'h644, 12'h544, 12'h543, 12'h544, 12'h544, 12'h533, 12'h433, 12'h433, 12'h323, 12'h332, 12'h333, 12'h323, 12'h433, 12'h333, 12'h222, 12'h444, 12'h333, 12'h323, 12'h323, 12'h333, 12'h323, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h333, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h545, 12'h455, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h444, 12'h545, 12'h454, 12'h555, 12'h545, 12'h555,
		12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h455, 12'h544, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h555, 12'h777, 12'h777, 12'h666, 12'h766, 12'h888, 12'h999, 12'h999, 12'h888, 12'h766, 12'h766, 12'h666, 12'h665, 12'h655, 12'h766, 12'h755, 12'h655, 12'h766, 12'h876, 12'h766, 12'h765, 12'h765, 12'h766, 12'h866, 12'h866, 12'h766, 12'h765, 12'h765, 12'h755, 12'h755, 12'h755, 12'h765, 12'h765, 12'h866, 12'h755, 12'h865, 12'h866, 12'h977, 12'h977, 12'h977, 12'h866, 12'h866, 12'h866, 12'h866, 12'h765, 12'h765, 12'h755, 12'h755, 12'h754, 12'h754, 12'h744, 12'h654, 12'h644, 12'h533, 12'h544, 12'h644, 12'h544, 12'h534, 12'h433, 12'h433, 12'h322, 12'h333, 12'h433, 12'h433, 12'h433, 12'h333, 12'h323, 12'h222, 12'h221, 12'h222, 12'h333, 12'h333, 12'h222, 12'h222, 12'h322, 12'h222, 12'h222, 12'h222, 12'h323, 12'h333, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h544, 12'h445, 12'h454, 12'h545, 12'h545,
		12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h544, 12'h444, 12'h444, 12'h455, 12'h544, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h544, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h445, 12'h545, 12'h665, 12'h666, 12'h777, 12'h877, 12'h989, 12'h989, 12'h878, 12'h888, 12'h766, 12'h655, 12'h665, 12'h665, 12'h766, 12'h766, 12'h755, 12'h655, 12'h755, 12'h765, 12'h755, 12'h756, 12'h766, 12'h866, 12'h866, 12'h866, 12'h865, 12'h866, 12'h966, 12'h976, 12'h966, 12'h866, 12'h976, 12'h966, 12'h966, 12'h976, 12'h966, 12'h866, 12'h966, 12'h966, 12'h976, 12'h866, 12'h866, 12'h865, 12'h865, 12'h865, 12'h855, 12'h755, 12'h755, 12'h855, 12'h755, 12'h754, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h322, 12'h222, 12'h211, 12'h322, 12'h333, 12'h323, 12'h222, 12'h333, 12'h433, 12'h223, 12'h222, 12'h323, 12'h333, 12'h444, 12'h445, 12'h555, 12'h455, 12'h555, 12'h455, 12'h455, 12'h555, 12'h555, 12'h455, 12'h445, 12'h555, 12'h455, 12'h545, 12'h555, 12'h444, 12'h445, 12'h445, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h545, 12'h545, 12'h455, 12'h445,
		12'h444, 12'h454, 12'h445, 12'h544, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h454, 12'h444, 12'h545, 12'h454, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h545, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h454, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h454, 12'h545, 12'h444, 12'h454, 12'h444, 12'h545, 12'h444, 12'h544, 12'h666, 12'h877, 12'h888, 12'h888, 12'h877, 12'h877, 12'h777, 12'h766, 12'h766, 12'h766, 12'h655, 12'h655, 12'h654, 12'h654, 12'h755, 12'h765, 12'h765, 12'h866, 12'h866, 12'h755, 12'h865, 12'h866, 12'h976, 12'h976, 12'h976, 12'h976, 12'h976, 12'hA76, 12'hA77, 12'h976, 12'hA76, 12'h976, 12'h966, 12'h976, 12'hA77, 12'h976, 12'h976, 12'h966, 12'h976, 12'h966, 12'hA76, 12'h976, 12'h966, 12'h966, 12'h966, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h755, 12'h755, 12'h744, 12'h744, 12'h744, 12'h644, 12'h644, 12'h755, 12'h644, 12'h533, 12'h644, 12'h644, 12'h533, 12'h433, 12'h433, 12'h433, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h323, 12'h222, 12'h333, 12'h444, 12'h333, 12'h222, 12'h333, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h445, 12'h454, 12'h555, 12'h445, 12'h454, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h445, 12'h555, 12'h444, 12'h454, 12'h555, 12'h444, 12'h455, 12'h455,
		12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h455, 12'h555, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h544, 12'h445, 12'h444, 12'h555, 12'h445, 12'h444, 12'h445, 12'h445, 12'h444, 12'h454, 12'h445, 12'h444, 12'h454, 12'h445, 12'h545, 12'h454, 12'h444, 12'h444, 12'h445, 12'h554, 12'h555, 12'h777, 12'h888, 12'h888, 12'h766, 12'h666, 12'h766, 12'h766, 12'h655, 12'h645, 12'h644, 12'h654, 12'h755, 12'h755, 12'h865, 12'h866, 12'h966, 12'h976, 12'h976, 12'h966, 12'h976, 12'h976, 12'hA76, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'hA77, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'h966, 12'h966, 12'h966, 12'h965, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h754, 12'h754, 12'h755, 12'h754, 12'h744, 12'h754, 12'h744, 12'h644, 12'h644, 12'h644, 12'h633, 12'h533, 12'h543, 12'h533, 12'h533, 12'h433, 12'h422, 12'h322, 12'h322, 12'h222, 12'h211, 12'h222, 12'h322, 12'h323, 12'h333, 12'h333, 12'h444, 12'h444, 12'h545, 12'h333, 12'h222, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h454, 12'h545, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h545, 12'h555, 12'h545, 12'h445, 12'h554, 12'h455, 12'h445, 12'h545,
		12'h444, 12'h445, 12'h544, 12'h454, 12'h445, 12'h444, 12'h444, 12'h555, 12'h454, 12'h444, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h544, 12'h445, 12'h444, 12'h455, 12'h444, 12'h454, 12'h445, 12'h544, 12'h454, 12'h445, 12'h454, 12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h554, 12'h445, 12'h444, 12'h545, 12'h555, 12'h555, 12'h545, 12'h555, 12'h767, 12'h989, 12'h888, 12'h877, 12'h766, 12'h666, 12'h545, 12'h655, 12'h544, 12'h544, 12'h654, 12'h754, 12'h865, 12'h876, 12'h976, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA87, 12'hA87, 12'hA87, 12'hA76, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA77, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h966, 12'h965, 12'h965, 12'h965, 12'h855, 12'h855, 12'h854, 12'h854, 12'h855, 12'h754, 12'h754, 12'h754, 12'h744, 12'h754, 12'h644, 12'h644, 12'h643, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h433, 12'h433, 12'h423, 12'h322, 12'h211, 12'h211, 12'h222, 12'h323, 12'h322, 12'h333, 12'h333, 12'h444, 12'h444, 12'h545, 12'h222, 12'h222, 12'h434, 12'h555, 12'h444, 12'h555, 12'h555, 12'h445, 12'h455, 12'h554, 12'h445, 12'h555, 12'h555, 12'h445, 12'h555, 12'h455, 12'h545, 12'h554, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h545, 12'h445, 12'h554, 12'h544,
		12'h444, 12'h444, 12'h445, 12'h544, 12'h454, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h454, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h445, 12'h444, 12'h454, 12'h444, 12'h545, 12'h444, 12'h455, 12'h544, 12'h445, 12'h454, 12'h545, 12'h444, 12'h554, 12'h445, 12'h444, 12'h454, 12'h445, 12'h445, 12'h554, 12'h445, 12'h454, 12'h555, 12'h445, 12'h444, 12'h555, 12'h777, 12'h777, 12'h888, 12'h878, 12'h777, 12'h766, 12'h656, 12'h544, 12'h655, 12'h655, 12'h655, 12'h866, 12'h976, 12'h987, 12'hA87, 12'hB98, 12'hA87, 12'hA87, 12'hA87, 12'hA77, 12'hA87, 12'hB87, 12'hA77, 12'hB87, 12'hB87, 12'hB87, 12'hA76, 12'hA76, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h965, 12'h965, 12'h855, 12'h854, 12'h855, 12'h854, 12'h854, 12'h755, 12'h754, 12'h754, 12'h754, 12'h754, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h643, 12'h533, 12'h533, 12'h533, 12'h433, 12'h423, 12'h322, 12'h312, 12'h222, 12'h222, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h444, 12'h444, 12'h333, 12'h333, 12'h444, 12'h555, 12'h555, 12'h544, 12'h444, 12'h555, 12'h555, 12'h445, 12'h555, 12'h454, 12'h444, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h455, 12'h555, 12'h554, 12'h555, 12'h554, 12'h455, 12'h545, 12'h554, 12'h454,
		12'h444, 12'h455, 12'h444, 12'h445, 12'h444, 12'h545, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h444, 12'h445, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h445, 12'h444, 12'h555, 12'h444, 12'h445, 12'h555, 12'h444, 12'h555, 12'h455, 12'h445, 12'h555, 12'h444, 12'h545, 12'h555, 12'h444, 12'h455, 12'h544, 12'h445, 12'h555, 12'h544, 12'h444, 12'h544, 12'h555, 12'h665, 12'h777, 12'h877, 12'h999, 12'h777, 12'h766, 12'h656, 12'h655, 12'h544, 12'h655, 12'h766, 12'h866, 12'hA88, 12'hA98, 12'hB98, 12'hB88, 12'hB98, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h965, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h755, 12'h754, 12'h855, 12'h754, 12'h754, 12'h754, 12'h744, 12'h643, 12'h644, 12'h644, 12'h644, 12'h633, 12'h533, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h322, 12'h212, 12'h222, 12'h221, 12'h222, 12'h322, 12'h222, 12'h222, 12'h333, 12'h555, 12'h444, 12'h333, 12'h334, 12'h555, 12'h444, 12'h445, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h555, 12'h545, 12'h454, 12'h555, 12'h545, 12'h455, 12'h545, 12'h544, 12'h455, 12'h545, 12'h444, 12'h454, 12'h555, 12'h444, 12'h444,
		12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h455, 12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h454, 12'h445, 12'h444, 12'h445, 12'h444, 12'h445, 12'h454, 12'h445, 12'h444, 12'h444, 12'h445, 12'h454, 12'h544, 12'h444, 12'h455, 12'h555, 12'h444, 12'h555, 12'h444, 12'h555, 12'h444, 12'h544, 12'h455, 12'h444, 12'h455, 12'h455, 12'h544, 12'h455, 12'h545, 12'h554, 12'h455, 12'h545, 12'h554, 12'h555, 12'h544, 12'h656, 12'h777, 12'h877, 12'h999, 12'h766, 12'h766, 12'h776, 12'h655, 12'h655, 12'h755, 12'h876, 12'h977, 12'h987, 12'hB98, 12'hB99, 12'hB98, 12'hB98, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hB87, 12'hA77, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hA76, 12'hA76, 12'hB77, 12'hA77, 12'hA86, 12'hB77, 12'hB87, 12'hB87, 12'hB87, 12'hA87, 12'hA87, 12'hA87, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA76, 12'h976, 12'h966, 12'h965, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h844, 12'h855, 12'h855, 12'h754, 12'h744, 12'h754, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h543, 12'h533, 12'h433, 12'h433, 12'h322, 12'h321, 12'h321, 12'h211, 12'h222, 12'h222, 12'h322, 12'h333, 12'h333, 12'h323, 12'h333, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h455, 12'h544, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h454, 12'h555, 12'h445, 12'h554, 12'h455, 12'h555, 12'h555, 12'h455, 12'h544, 12'h454, 12'h454,
		12'h445, 12'h444, 12'h454, 12'h545, 12'h444, 12'h455, 12'h544, 12'h444, 12'h455, 12'h444, 12'h544, 12'h445, 12'h554, 12'h444, 12'h454, 12'h545, 12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h455, 12'h445, 12'h444, 12'h445, 12'h554, 12'h445, 12'h445, 12'h554, 12'h455, 12'h445, 12'h555, 12'h555, 12'h444, 12'h545, 12'h555, 12'h444, 12'h455, 12'h545, 12'h455, 12'h545, 12'h554, 12'h445, 12'h555, 12'h555, 12'h555, 12'h766, 12'h777, 12'h766, 12'h766, 12'h766, 12'h887, 12'h555, 12'h766, 12'h877, 12'h877, 12'hA88, 12'hA98, 12'hB99, 12'hCA9, 12'hCA9, 12'hB99, 12'hC99, 12'hC98, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB88, 12'hB87, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA87, 12'hB87, 12'hB87, 12'hA77, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA87, 12'hA87, 12'hA77, 12'hA76, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h855, 12'h754, 12'h855, 12'h754, 12'h754, 12'h754, 12'h754, 12'h744, 12'h744, 12'h644, 12'h643, 12'h643, 12'h644, 12'h543, 12'h533, 12'h533, 12'h433, 12'h432, 12'h422, 12'h322, 12'h322, 12'h322, 12'h222, 12'h322, 12'h333, 12'h444, 12'h433, 12'h333, 12'h444, 12'h333, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h454, 12'h555, 12'h545, 12'h454, 12'h555, 12'h555,
		12'h445, 12'h444, 12'h455, 12'h444, 12'h445, 12'h554, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h444, 12'h445, 12'h444, 12'h444, 12'h555, 12'h444, 12'h444, 12'h445, 12'h554, 12'h444, 12'h545, 12'h554, 12'h445, 12'h454, 12'h545, 12'h454, 12'h545, 12'h555, 12'h454, 12'h545, 12'h555, 12'h454, 12'h445, 12'h555, 12'h554, 12'h445, 12'h545, 12'h555, 12'h455, 12'h444, 12'h545, 12'h555, 12'h545, 12'h555, 12'h666, 12'h666, 12'h777, 12'h878, 12'h766, 12'h877, 12'h767, 12'h988, 12'h988, 12'h987, 12'hA98, 12'hB99, 12'hBA9, 12'hCA9, 12'hCAA, 12'hCA9, 12'hCA9, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA87, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h965, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h755, 12'h855, 12'h855, 12'h855, 12'h754, 12'h744, 12'h754, 12'h744, 12'h644, 12'h643, 12'h644, 12'h644, 12'h544, 12'h543, 12'h533, 12'h433, 12'h433, 12'h433, 12'h333, 12'h322, 12'h333, 12'h333, 12'h323, 12'h444, 12'h544, 12'h334, 12'h333, 12'h333, 12'h111, 12'h333, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h545, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h554, 12'h545, 12'h555, 12'h455, 12'h544, 12'h555, 12'h455, 12'h545, 12'h554, 12'h555, 12'h455, 12'h554, 12'h555, 12'h445, 12'h555, 12'h455, 12'h545, 12'h455, 12'h555, 12'h444, 12'h445, 12'h454, 12'h545, 12'h454, 12'h545, 12'h455, 12'h555, 12'h444, 12'h555, 12'h445, 12'h555, 12'h545, 12'h454, 12'h555, 12'h555, 12'h455, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h766, 12'h877, 12'h777, 12'h777, 12'h988, 12'h988, 12'h988, 12'h988, 12'hA99, 12'hBA9, 12'hCAA, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB88, 12'hB87, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'hA76, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h965, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h855, 12'h854, 12'h754, 12'h744, 12'h744, 12'h644, 12'h644, 12'h633, 12'h643, 12'h644, 12'h644, 12'h543, 12'h533, 12'h433, 12'h433, 12'h433, 12'h322, 12'h322, 12'h222, 12'h322, 12'h333, 12'h444, 12'h444, 12'h222, 12'h223, 12'h222, 12'h222, 12'h444, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h455, 12'h545, 12'h454, 12'h555, 12'h545, 12'h455, 12'h555, 12'h455, 12'h555, 12'h545, 12'h454, 12'h555, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h554, 12'h455, 12'h545, 12'h455, 12'h455, 12'h545, 12'h555, 12'h455, 12'h545, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h545, 12'h555, 12'h555, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h777, 12'h999, 12'h766, 12'h877, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'hA98, 12'hB99, 12'hBA9, 12'hCAA, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hC99, 12'hCA8, 12'hCA9, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hB98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC88, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hC88, 12'hB98, 12'hB98, 12'hB98, 12'hB98, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB77, 12'hA77, 12'hA77, 12'hA77, 12'hA66, 12'h966, 12'h966, 12'h966, 12'h965, 12'h965, 12'h955, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h754, 12'h755, 12'h744, 12'h744, 12'h744, 12'h644, 12'h643, 12'h643, 12'h644, 12'h644, 12'h533, 12'h533, 12'h432, 12'h433, 12'h423, 12'h322, 12'h322, 12'h322, 12'h333, 12'h333, 12'h333, 12'h222, 12'h222, 12'h223, 12'h122, 12'h333, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h455, 12'h545, 12'h455, 12'h555, 12'h555, 12'h445, 12'h554, 12'h445, 12'h455, 12'h545, 12'h445, 12'h455, 12'h545, 12'h454, 12'h555, 12'h445, 12'h445, 12'h554, 12'h545, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h655, 12'h766, 12'h878, 12'h777, 12'h877, 12'h988, 12'hA99, 12'hBAA, 12'hBA9, 12'hBA9, 12'hBAA, 12'hBAA, 12'hBA9, 12'hBA9, 12'hCAA, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hDA9, 12'hD99, 12'hC99, 12'hCA9, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC88, 12'hB88, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC99, 12'hC98, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hA77, 12'hA76, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h966, 12'h965, 12'h965, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h854, 12'h744, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h433, 12'h433, 12'h323, 12'h333, 12'h323, 12'h322, 12'h323, 12'h333, 12'h222, 12'h222, 12'h222, 12'h112, 12'h222, 12'h444, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h545, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h455, 12'h545, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h545, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h666, 12'h665, 12'h666, 12'h666, 12'h877, 12'h888, 12'h988, 12'hA99, 12'hAAA, 12'hAAA, 12'hBAA, 12'hBAA, 12'hCAA, 12'hCBA, 12'hCAA, 12'hCAA, 12'hCA9, 12'hCA9, 12'hCA9, 12'hDA9, 12'hCA9, 12'hDA9, 12'hC98, 12'hDA9, 12'hDA9, 12'hC99, 12'hC99, 12'hCA9, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB88, 12'hB77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h966, 12'h966, 12'h965, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h854, 12'h754, 12'h744, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h643, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h322, 12'h433, 12'h333, 12'h222, 12'h223, 12'h222, 12'h222, 12'h122, 12'h333, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h566, 12'h555, 12'h565, 12'h566, 12'h666, 12'h666, 12'h676, 12'h888, 12'h888, 12'h988, 12'hAAA, 12'hAAA, 12'hBAA, 12'hBAA, 12'hCBB, 12'hCBB, 12'hCBA, 12'hCAA, 12'hCA9, 12'hDA9, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hC99, 12'hC99, 12'hCA9, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hCA9, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC89, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h966, 12'h966, 12'h966, 12'h966, 12'h965, 12'h955, 12'h855, 12'h855, 12'h855, 12'h754, 12'h754, 12'h754, 12'h754, 12'h754, 12'h744, 12'h644, 12'h643, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h222, 12'h222, 12'h111, 12'h111, 12'h222, 12'h223, 12'h444, 12'h555, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h998, 12'h999, 12'hAAA, 12'hBBA, 12'hCBB, 12'hCBB, 12'hCBB, 12'hDBB, 12'hCBA, 12'hCBA, 12'hCA9, 12'hDAA, 12'hDA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hDA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hD99, 12'hCA9, 12'hDA9, 12'hD99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB77, 12'hA77, 12'hA76, 12'hA66, 12'hA66, 12'hA76, 12'hA66, 12'hA76, 12'h966, 12'h966, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h854, 12'h854, 12'h744, 12'h754, 12'h754, 12'h744, 12'h644, 12'h644, 12'h543, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h323, 12'h222, 12'h112, 12'h111, 12'h212, 12'h333, 12'h444, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h566, 12'h566, 12'h566, 12'h566, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h778, 12'h999, 12'hA99, 12'hA99, 12'hBBA, 12'hCBB, 12'hDCC, 12'hCBB, 12'hCBB, 12'hDBB, 12'hDBA, 12'hCBA, 12'hCAA, 12'hDBA, 12'hDB9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hCAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hD99, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hC99, 12'hC99, 12'hD99, 12'hC99, 12'hC99, 12'hD99, 12'hC99, 12'hD99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC98, 12'hC88, 12'hB88, 12'hB88, 12'hB87, 12'hB77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA66, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h965, 12'h855, 12'h855, 12'h855, 12'h854, 12'h854, 12'h854, 12'h854, 12'h754, 12'h744, 12'h744, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h433, 12'h223, 12'h222, 12'h111, 12'h222, 12'h444, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h556, 12'h566, 12'h556, 12'h566, 12'h556, 12'h555, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h565, 12'h556, 12'h566, 12'h566, 12'h656, 12'h565, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h777, 12'h898, 12'hAA9, 12'hCBB, 12'hCBB, 12'hCCC, 12'hCBB, 12'hCBB, 12'hCBA, 12'hDBB, 12'hDBB, 12'hDBA, 12'hCBA, 12'hCA9, 12'hDAA, 12'hDBA, 12'hDB9, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hDA9, 12'hD9A, 12'hCA9, 12'hCA9, 12'hD99, 12'hDA9, 12'hC99, 12'hD99, 12'hD99, 12'hC99, 12'hD99, 12'hD99, 12'hC99, 12'hDA9, 12'hC99, 12'hD99, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hB88, 12'hB88, 12'hB87, 12'hB77, 12'hB77, 12'hA77, 12'hA76, 12'hA76, 12'h966, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h854, 12'h754, 12'h754, 12'h744, 12'h644, 12'h644, 12'h543, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h443, 12'h444, 12'h544, 12'h444, 12'h223, 12'h222, 12'h111, 12'h222, 12'h444, 12'h666, 12'h556, 12'h555, 12'h666, 12'h666, 12'h555, 12'h555, 12'h566, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555,
		12'h555, 12'h555, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h656, 12'h655, 12'h566, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h566, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'hBBB, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCCC, 12'hCBB, 12'hCBB, 12'hDCB, 12'hDBB, 12'hDBA, 12'hCAA, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDA9, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hCA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hC99, 12'hC99, 12'hCA9, 12'hD99, 12'hDAA, 12'hDA9, 12'hDA9, 12'hC99, 12'hCA9, 12'hDA9, 12'hDA9, 12'hC99, 12'hDA9, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hB88, 12'hB77, 12'hA77, 12'hA66, 12'hA66, 12'hA77, 12'hA77, 12'h966, 12'h966, 12'h966, 12'h966, 12'h965, 12'h855, 12'h855, 12'h855, 12'h865, 12'h865, 12'h955, 12'h855, 12'h854, 12'h754, 12'h744, 12'h644, 12'h643, 12'h534, 12'h533, 12'h533, 12'h433, 12'h433, 12'h544, 12'h544, 12'h544, 12'h545, 12'h444, 12'h433, 12'h212, 12'h222, 12'h222, 12'h445, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h655, 12'h655, 12'h666, 12'h655, 12'h555, 12'h656, 12'h555, 12'h555,
		12'h556, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h556, 12'h555, 12'h555, 12'h556, 12'h566, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h777, 12'h999, 12'hBAA, 12'hCBB, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hCBB, 12'hDBB, 12'hDCB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hDBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hC99, 12'hD99, 12'hC99, 12'hDA9, 12'hD99, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hC98, 12'hC99, 12'hD99, 12'hDA9, 12'hC99, 12'hC98, 12'hC98, 12'hC88, 12'hB77, 12'hA77, 12'hA76, 12'hA77, 12'hA77, 12'hA77, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h965, 12'h865, 12'h855, 12'h855, 12'h865, 12'h965, 12'h855, 12'h855, 12'h855, 12'h754, 12'h744, 12'h644, 12'h644, 12'h543, 12'h533, 12'h533, 12'h433, 12'h533, 12'h534, 12'h544, 12'h544, 12'h545, 12'h544, 12'h333, 12'h323, 12'h222, 12'h222, 12'h445, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h666, 12'h666, 12'h656, 12'h556, 12'h566, 12'h656, 12'h555, 12'h566, 12'h655, 12'h556, 12'h665, 12'h655, 12'h555, 12'h555,
		12'h565, 12'h556, 12'h665, 12'h565, 12'h566, 12'h666, 12'h555, 12'h566, 12'h555, 12'h665, 12'h566, 12'h656, 12'h565, 12'h666, 12'h666, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h677, 12'h777, 12'h777, 12'h999, 12'hBBB, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hDCC, 12'hDBB, 12'hDBB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hCAA, 12'hD99, 12'hD99, 12'hC99, 12'hD99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hD99, 12'hCA9, 12'hC99, 12'hD99, 12'hC98, 12'hC98, 12'hC99, 12'hC99, 12'hD99, 12'hC99, 12'hC99, 12'hC88, 12'hB87, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB87, 12'hA76, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h965, 12'h855, 12'h855, 12'h965, 12'h965, 12'h855, 12'h855, 12'h854, 12'h855, 12'h754, 12'h644, 12'h644, 12'h643, 12'h533, 12'h533, 12'h533, 12'h433, 12'h543, 12'h444, 12'h544, 12'h544, 12'h545, 12'h333, 12'h333, 12'h323, 12'h222, 12'h444, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h566, 12'h656, 12'h655, 12'h666, 12'h656, 12'h655, 12'h566, 12'h656, 12'h655, 12'h665,
		12'h555, 12'h656, 12'h556, 12'h555, 12'h655, 12'h556, 12'h565, 12'h656, 12'h556, 12'h555, 12'h666, 12'h556, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h677, 12'h677, 12'h667, 12'h677, 12'h677, 12'h677, 12'h666, 12'h777, 12'h666, 12'h888, 12'hBBB, 12'hCCC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hDBC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDBB, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEAA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hDBB, 12'hEBB, 12'hEBB, 12'hDBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hCA9, 12'hC99, 12'hD99, 12'hDA9, 12'hC99, 12'hD99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hC99, 12'hC99, 12'hDA9, 12'hC99, 12'hC99, 12'hC98, 12'hC88, 12'hB87, 12'hA77, 12'hB87, 12'hB77, 12'hB87, 12'hA77, 12'hA76, 12'hA76, 12'h966, 12'h965, 12'h966, 12'h965, 12'h855, 12'h955, 12'h965, 12'h855, 12'h854, 12'h855, 12'h854, 12'h744, 12'h644, 12'h644, 12'h644, 12'h533, 12'h544, 12'h433, 12'h533, 12'h544, 12'h544, 12'h544, 12'h444, 12'h545, 12'h444, 12'h434, 12'h333, 12'h323, 12'h444, 12'h666, 12'h667, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h565, 12'h666, 12'h655, 12'h666, 12'h655, 12'h656, 12'h666,
		12'h666, 12'h566, 12'h566, 12'h656, 12'h665, 12'h566, 12'h656, 12'h666, 12'h666, 12'h666, 12'h665, 12'h566, 12'h655, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h666, 12'h667, 12'h667, 12'h666, 12'h666, 12'h667, 12'h676, 12'h676, 12'h676, 12'h666, 12'h677, 12'h677, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'hAAA, 12'hBBB, 12'hCCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCB, 12'hDCB, 12'hDBB, 12'hEBA, 12'hDBB, 12'hDBA, 12'hEBB, 12'hDBA, 12'hDBB, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBB, 12'hEBB, 12'hECB, 12'hDBB, 12'hECB, 12'hECB, 12'hDBA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBA, 12'hDAA, 12'hDAB, 12'hDBB, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC99, 12'hD99, 12'hD99, 12'hDA9, 12'hDAA, 12'hD99, 12'hD99, 12'hC99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC99, 12'hC99, 12'hC99, 12'hD99, 12'hDA9, 12'hDA9, 12'hD99, 12'hC98, 12'hC88, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB88, 12'hA77, 12'hA77, 12'hA76, 12'h966, 12'h966, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h755, 12'h754, 12'h644, 12'h643, 12'h633, 12'h533, 12'h433, 12'h543, 12'h433, 12'h433, 12'h433, 12'h534, 12'h544, 12'h444, 12'h444, 12'h433, 12'h333, 12'h333, 12'h444, 12'h666, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h556, 12'h666, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666,
		12'h556, 12'h665, 12'h565, 12'h656, 12'h566, 12'h565, 12'h656, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h676, 12'h777, 12'h667, 12'h677, 12'h676, 12'h677, 12'h667, 12'h677, 12'h677, 12'h677, 12'h776, 12'h777, 12'h677, 12'h776, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'hBAB, 12'hCBC, 12'hCCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hDCC, 12'hECB, 12'hDBB, 12'hDBA, 12'hEBB, 12'hEBB, 12'hDBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBB, 12'hECB, 12'hECC, 12'hECC, 12'hECB, 12'hEBB, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hCA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hCA9, 12'hD9A, 12'hC99, 12'hC99, 12'hD99, 12'hDAA, 12'hDAA, 12'hEAA, 12'hDA9, 12'hDA9, 12'hC99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDA9, 12'hC99, 12'hC98, 12'hC88, 12'hB88, 12'hB87, 12'hB87, 12'hB88, 12'hB88, 12'hB77, 12'hA77, 12'hA77, 12'hA77, 12'h966, 12'h966, 12'h965, 12'h965, 12'h865, 12'h865, 12'h865, 12'h855, 12'h855, 12'h755, 12'h754, 12'h644, 12'h644, 12'h543, 12'h533, 12'h533, 12'h544, 12'h433, 12'h533, 12'h433, 12'h433, 12'h533, 12'h434, 12'h444, 12'h444, 12'h333, 12'h333, 12'h555, 12'h666, 12'h777, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h656, 12'h666, 12'h666, 12'h656, 12'h666, 12'h666, 12'h666,
		12'h666, 12'h656, 12'h556, 12'h666, 12'h656, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h666, 12'h776, 12'h767, 12'h777, 12'h776, 12'h777, 12'h676, 12'h676, 12'h767, 12'h767, 12'h677, 12'h777, 12'h767, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'hBBB, 12'hCCC, 12'hCCC, 12'hDDD, 12'hEDD, 12'hECC, 12'hDCB, 12'hDBB, 12'hDBB, 12'hECB, 12'hEBA, 12'hEBB, 12'hDBB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hECB, 12'hECC, 12'hECB, 12'hDBB, 12'hC99, 12'hB99, 12'hB98, 12'hB88, 12'hB98, 12'hB99, 12'hCA9, 12'hCA9, 12'hB99, 12'hB98, 12'hB88, 12'hB88, 12'hB99, 12'hC99, 12'hDAA, 12'hCAA, 12'hCA9, 12'hDAA, 12'hDAB, 12'hDAA, 12'hDAA, 12'hDAA, 12'hC9A, 12'hDAA, 12'hC99, 12'hCA9, 12'hDA9, 12'hEBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hC99, 12'hC88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB77, 12'hA77, 12'hA77, 12'hA76, 12'h966, 12'h966, 12'h966, 12'h966, 12'h866, 12'h855, 12'h855, 12'h865, 12'h755, 12'h755, 12'h754, 12'h644, 12'h634, 12'h544, 12'h543, 12'h533, 12'h544, 12'h533, 12'h534, 12'h533, 12'h443, 12'h433, 12'h544, 12'h434, 12'h444, 12'h444, 12'h333, 12'h555, 12'h777, 12'h777, 12'h666, 12'h677, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h656, 12'h666, 12'h665, 12'h666, 12'h666,
		12'h566, 12'h555, 12'h666, 12'h566, 12'h656, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h666, 12'h667, 12'h667, 12'h667, 12'h666, 12'h667, 12'h777, 12'h777, 12'h667, 12'h677, 12'h767, 12'h767, 12'h677, 12'h767, 12'h776, 12'h777, 12'h676, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'hBBB, 12'hCCC, 12'hCCC, 12'hEDD, 12'hDDD, 12'hDCC, 12'hECC, 12'hDCB, 12'hDBB, 12'hDBA, 12'hEBA, 12'hDBB, 12'hEBA, 12'hECB, 12'hDBB, 12'hECB, 12'hDBB, 12'hDBB, 12'hECB, 12'hECB, 12'hDBB, 12'hDBA, 12'hCAA, 12'hCAA, 12'hCA9, 12'hB99, 12'hB98, 12'hB98, 12'hB99, 12'hB88, 12'hA88, 12'hA88, 12'hB88, 12'hB88, 12'hA88, 12'hA77, 12'hA77, 12'hB88, 12'hB89, 12'hB88, 12'hC99, 12'hDAA, 12'hCAA, 12'hDAA, 12'hDAA, 12'hCAA, 12'hCAA, 12'hC99, 12'hDAA, 12'hDAA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDA9, 12'hCA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hC98, 12'hC98, 12'hC88, 12'hB88, 12'hB88, 12'hB87, 12'hA77, 12'hA77, 12'h977, 12'h966, 12'h855, 12'h866, 12'h855, 12'h755, 12'h755, 12'h755, 12'h755, 12'h755, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h533, 12'h443, 12'h543, 12'h544, 12'h534, 12'h433, 12'h544, 12'h433, 12'h444, 12'h444, 12'h433, 12'h444, 12'h334, 12'h555, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h777, 12'h777, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666,
		12'h556, 12'h665, 12'h665, 12'h566, 12'h666, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h776, 12'h677, 12'h677, 12'h776, 12'h677, 12'h667, 12'h666, 12'h777, 12'h667, 12'h776, 12'h677, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'hBBB, 12'hCCC, 12'hDCC, 12'hEDD, 12'hEDC, 12'hECC, 12'hECC, 12'hECB, 12'hDBB, 12'hEBA, 12'hDBB, 12'hEBB, 12'hECB, 12'hEBB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hCAA, 12'hCAA, 12'hDAA, 12'hCA9, 12'hC99, 12'hC99, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hA78, 12'hB88, 12'hB88, 12'hB89, 12'hB88, 12'hC99, 12'hC99, 12'hC99, 12'hC9A, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDBA, 12'hEBB, 12'hDBA, 12'hDAA, 12'hDAA, 12'hC99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hC88, 12'hB88, 12'hB77, 12'hB77, 12'hA77, 12'h966, 12'h966, 12'h865, 12'h855, 12'h755, 12'h744, 12'h744, 12'h744, 12'h754, 12'h755, 12'h755, 12'h744, 12'h645, 12'h644, 12'h533, 12'h533, 12'h534, 12'h544, 12'h533, 12'h533, 12'h533, 12'h544, 12'h544, 12'h533, 12'h433, 12'h433, 12'h534, 12'h433, 12'h444, 12'h444, 12'h444, 12'h444, 12'h666, 12'h777, 12'h666, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h776, 12'h767, 12'h666, 12'h666, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666,
		12'h666, 12'h666, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h767, 12'h676, 12'h767, 12'h666, 12'h776, 12'h767, 12'h677, 12'h776, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'h999, 12'hCBB, 12'hDCC, 12'hDDD, 12'hEDD, 12'hEDD, 12'hECC, 12'hECC, 12'hECB, 12'hECB, 12'hEBB, 12'hECA, 12'hECB, 12'hDBB, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hDBB, 12'hDBA, 12'hDBB, 12'hDBB, 12'hDBB, 12'hDAA, 12'hDAA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC99, 12'hC88, 12'hC88, 12'hC88, 12'hB88, 12'hB88, 12'hC88, 12'hC99, 12'hC88, 12'hC88, 12'hC99, 12'hC99, 12'hC99, 12'hD99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hC99, 12'hC99, 12'hC99, 12'hCA9, 12'hDA9, 12'hD99, 12'hC98, 12'hB88, 12'hB87, 12'hA77, 12'hA77, 12'h966, 12'h855, 12'h855, 12'h744, 12'h744, 12'h644, 12'h533, 12'h533, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h534, 12'h544, 12'h533, 12'h533, 12'h433, 12'h433, 12'h543, 12'h544, 12'h533, 12'h433, 12'h433, 12'h443, 12'h444, 12'h545, 12'h444, 12'h444, 12'h444, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h777, 12'h777, 12'h777, 12'h766, 12'h766, 12'h766, 12'h666, 12'h666, 12'h766, 12'h666, 12'h666,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h676, 12'h767, 12'h667, 12'h677, 12'h667, 12'h766, 12'h677, 12'h666, 12'h777, 12'h777, 12'h667, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'hA99, 12'hCCC, 12'hDDD, 12'hEDD, 12'hEDD, 12'hEDD, 12'hEDC, 12'hECC, 12'hECB, 12'hECB, 12'hEBB, 12'hEBA, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hECC, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBB, 12'hDBB, 12'hDBB, 12'hEBB, 12'hDBB, 12'hDBB, 12'hDBB, 12'hDBA, 12'hEBA, 12'hDAA, 12'hDAA, 12'hD99, 12'hC99, 12'hC99, 12'hC89, 12'hD99, 12'hC99, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hC99, 12'hD99, 12'hDA9, 12'hD99, 12'hDAA, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hC98, 12'hC88, 12'hC98, 12'hC99, 12'hC99, 12'hC88, 12'hB87, 12'hB77, 12'hA66, 12'h966, 12'h855, 12'h855, 12'h744, 12'h644, 12'h644, 12'h644, 12'h633, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h533, 12'h534, 12'h544, 12'h544, 12'h533, 12'h433, 12'h443, 12'h533, 12'h544, 12'h534, 12'h533, 12'h433, 12'h433, 12'h544, 12'h555, 12'h444, 12'h444, 12'h444, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h676, 12'h777, 12'h767, 12'h767, 12'h766, 12'h767, 12'h766, 12'h766, 12'h666, 12'h666,
		12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h766, 12'h777, 12'h677, 12'h776, 12'h777, 12'h667, 12'h777, 12'h777, 12'h676, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h877, 12'hA99, 12'hDBB, 12'hDCC, 12'hDCB, 12'hCAA, 12'hA88, 12'h987, 12'h876, 12'hBA9, 12'hDCC, 12'hDDD, 12'hEEE, 12'hEDD, 12'hEDD, 12'hEDD, 12'hECC, 12'hECB, 12'hECB, 12'hECB, 12'hDBB, 12'hDBB, 12'hEBB, 12'hECB, 12'hECB, 12'hEBB, 12'hDBB, 12'hDBB, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hEBA, 12'hDAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hD99, 12'hD99, 12'hC98, 12'hC88, 12'hC87, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC98, 12'hC99, 12'hC98, 12'hC98, 12'hC98, 12'hC99, 12'hD99, 12'hDA9, 12'hD99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hEBA, 12'hEAA, 12'hEAA, 12'hDA9, 12'hB88, 12'hB87, 12'hB88, 12'hC88, 12'hC88, 12'hB88, 12'hB77, 12'hA67, 12'h965, 12'h754, 12'h744, 12'h643, 12'h643, 12'h633, 12'h644, 12'h744, 12'h744, 12'h855, 12'h855, 12'h966, 12'h967, 12'h966, 12'h966, 12'h866, 12'h755, 12'h755, 12'h644, 12'h644, 12'h544, 12'h544, 12'h533, 12'h433, 12'h433, 12'h533, 12'h443, 12'h433, 12'h433, 12'h433, 12'h544, 12'h544, 12'h544, 12'h444, 12'h555, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h677, 12'h777, 12'h767, 12'h766, 12'h666, 12'h766, 12'h766,
		12'h666, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h666, 12'h777, 12'h777, 12'h767, 12'h677, 12'h777, 12'h777, 12'h767, 12'h667, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h878, 12'h777, 12'h767, 12'hA88, 12'hDBB, 12'hDBA, 12'hDA9, 12'hD99, 12'hD99, 12'hEAA, 12'hEAA, 12'hDA9, 12'hC99, 12'hCAA, 12'hCCB, 12'hDDC, 12'hEED, 12'hEEE, 12'hEDD, 12'hEDD, 12'hECC, 12'hECC, 12'hECB, 12'hECB, 12'hEBB, 12'hDCB, 12'hECB, 12'hECC, 12'hECB, 12'hEBB, 12'hDBA, 12'hDBB, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hEBA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC98, 12'hC98, 12'hD98, 12'hC98, 12'hC87, 12'hC88, 12'hC88, 12'hC88, 12'hB87, 12'hB87, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC89, 12'hD99, 12'hD99, 12'hC99, 12'hD99, 12'hDA9, 12'hDAA, 12'hDBA, 12'hDAA, 12'hEAA, 12'hDA9, 12'hD99, 12'hB77, 12'hB77, 12'hB77, 12'hA77, 12'hA77, 12'hA76, 12'h966, 12'h855, 12'h744, 12'h633, 12'h633, 12'h532, 12'h633, 12'h633, 12'h744, 12'h955, 12'hA76, 12'hA66, 12'hA76, 12'hA77, 12'hB77, 12'hA77, 12'hA66, 12'h966, 12'h866, 12'h855, 12'h755, 12'h654, 12'h644, 12'h544, 12'h543, 12'h433, 12'h433, 12'h433, 12'h534, 12'h433, 12'h433, 12'h433, 12'h544, 12'h555, 12'h544, 12'h444, 12'h655, 12'h777, 12'h777, 12'h877, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h766,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h666, 12'h777, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h878, 12'h877, 12'h877, 12'hA88, 12'hDAA, 12'hD99, 12'hB67, 12'hA66, 12'hB77, 12'hC88, 12'hD88, 12'hE99, 12'hEBA, 12'hDAA, 12'hCAA, 12'hEDC, 12'hFEE, 12'hEED, 12'hEEE, 12'hEDD, 12'hEDD, 12'hEDD, 12'hECC, 12'hECB, 12'hECB, 12'hECC, 12'hECC, 12'hECB, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDBA, 12'hDAA, 12'hD99, 12'hDAA, 12'hC99, 12'hC89, 12'hC88, 12'hC88, 12'hB77, 12'h966, 12'hA66, 12'hA66, 12'hB77, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hD98, 12'hC98, 12'hD99, 12'hDAA, 12'hDAA, 12'hEAA, 12'hEBA, 12'hDAA, 12'hDA9, 12'hC98, 12'hB77, 12'hA66, 12'h965, 12'h965, 12'h966, 12'h855, 12'h855, 12'h744, 12'h533, 12'h522, 12'h532, 12'h744, 12'h855, 12'h966, 12'hA76, 12'hA77, 12'hB77, 12'hB77, 12'hB87, 12'hB88, 12'hB87, 12'hA77, 12'hA77, 12'h966, 12'h865, 12'h855, 12'h755, 12'h754, 12'h644, 12'h544, 12'h543, 12'h433, 12'h433, 12'h533, 12'h534, 12'h433, 12'h534, 12'h433, 12'h544, 12'h555, 12'h545, 12'h444, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h666, 12'h777, 12'h666, 12'h777, 12'h777, 12'h677, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h877, 12'h977, 12'hC99, 12'hD99, 12'hB67, 12'hD77, 12'hE88, 12'hE99, 12'hD98, 12'hD88, 12'hD88, 12'hC98, 12'hD99, 12'hDBA, 12'hECB, 12'hEDD, 12'hEDD, 12'hFED, 12'hDCC, 12'hDCC, 12'hECC, 12'hECB, 12'hECB, 12'hECC, 12'hECC, 12'hECC, 12'hECC, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hCA9, 12'hC99, 12'hDA9, 12'hC99, 12'hB88, 12'hB77, 12'hA77, 12'h966, 12'h845, 12'h745, 12'h745, 12'h745, 12'h745, 12'h745, 12'h966, 12'h855, 12'h855, 12'h966, 12'hA77, 12'hB77, 12'hB88, 12'hB77, 12'hC87, 12'hC88, 12'hC88, 12'hD98, 12'hD98, 12'hD99, 12'hDAA, 12'hEAA, 12'hEBA, 12'hDBA, 12'hEAA, 12'hDA9, 12'hC99, 12'hB77, 12'h965, 12'h854, 12'h744, 12'h633, 12'h633, 12'h634, 12'h533, 12'h523, 12'h644, 12'h755, 12'h855, 12'h966, 12'hA77, 12'hA77, 12'hB77, 12'hB88, 12'hB88, 12'hB88, 12'hB77, 12'hA77, 12'hA77, 12'hA66, 12'h966, 12'h855, 12'h855, 12'h755, 12'h644, 12'h633, 12'h533, 12'h544, 12'h533, 12'h433, 12'h433, 12'h543, 12'h433, 12'h433, 12'h433, 12'h544, 12'h655, 12'h444, 12'h433, 12'h777, 12'h788, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h666, 12'h667, 12'h666, 12'h777, 12'h667, 12'h676, 12'h777, 12'h777, 12'h767, 12'h776, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h787, 12'h887, 12'h776, 12'h876, 12'hC99, 12'hD88, 12'hD88, 12'hD88, 12'hE99, 12'hE99, 12'hE99, 12'hEA9, 12'hDA9, 12'hD99, 12'hC88, 12'hDA9, 12'hDBA, 12'hECB, 12'hECC, 12'hECC, 12'hDBB, 12'hDBB, 12'hECB, 12'hECB, 12'hDCB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hDBB, 12'hEBA, 12'hDAA, 12'hDA9, 12'hCA9, 12'hC99, 12'hC98, 12'hB87, 12'hA66, 12'hA66, 12'hA66, 12'h855, 12'h866, 12'hA78, 12'h755, 12'h867, 12'h544, 12'h655, 12'h544, 12'h655, 12'h755, 12'h856, 12'h855, 12'h855, 12'h955, 12'h956, 12'hA77, 12'hB66, 12'hB76, 12'hB77, 12'hC87, 12'hD98, 12'hD99, 12'hD99, 12'hDA9, 12'hEAA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDA9, 12'hC98, 12'hA76, 12'h855, 12'h743, 12'h633, 12'h532, 12'h533, 12'h523, 12'h423, 12'h533, 12'h745, 12'h855, 12'h755, 12'h744, 12'h744, 12'h855, 12'h966, 12'h976, 12'hA77, 12'hA88, 12'hA78, 12'hA77, 12'hA77, 12'h966, 12'h856, 12'h855, 12'h855, 12'h745, 12'h644, 12'h643, 12'h644, 12'h533, 12'h433, 12'h433, 12'h533, 12'h534, 12'h544, 12'h433, 12'h433, 12'h544, 12'h655, 12'h444, 12'h433, 12'h777, 12'h787, 12'h888, 12'h777, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h666, 12'h666, 12'h667, 12'h667, 12'h666, 12'h667, 12'h667, 12'h666, 12'h767, 12'h777, 12'h676, 12'h767, 12'h767, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h778, 12'h777, 12'h887, 12'h877, 12'h876, 12'hDAA, 12'hD99, 12'hC88, 12'hD88, 12'hE99, 12'hE99, 12'hD99, 12'hDA9, 12'hEBA, 12'hEAA, 12'hE99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hECB, 12'hECC, 12'hECB, 12'hECB, 12'hECC, 12'hECC, 12'hECB, 12'hEBB, 12'hDAA, 12'hEBA, 12'hDBA, 12'hEBA, 12'hDAA, 12'hC99, 12'hB88, 12'hB87, 12'hA76, 12'h965, 12'h955, 12'h844, 12'h966, 12'hCAA, 12'hDBB, 12'h866, 12'hCAB, 12'h877, 12'h323, 12'h322, 12'h666, 12'h744, 12'hA77, 12'hB88, 12'h966, 12'h955, 12'h955, 12'hA66, 12'hB66, 12'hB77, 12'hB77, 12'hC87, 12'hD99, 12'hDA9, 12'hD99, 12'hEAA, 12'hEBA, 12'hDAA, 12'hEAA, 12'hDAA, 12'hD99, 12'hC88, 12'hA66, 12'h844, 12'h633, 12'h522, 12'h533, 12'h422, 12'h422, 12'h433, 12'h633, 12'h633, 12'h533, 12'h633, 12'h866, 12'h866, 12'h866, 12'h755, 12'h643, 12'h644, 12'h534, 12'h533, 12'h645, 12'h744, 12'h644, 12'h745, 12'h755, 12'h745, 12'h644, 12'h533, 12'h533, 12'h533, 12'h433, 12'h533, 12'h533, 12'h534, 12'h534, 12'h543, 12'h433, 12'h534, 12'h544, 12'h544, 12'h333, 12'h333, 12'h777, 12'h888, 12'h778, 12'h777, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h666, 12'h667, 12'h666, 12'h666, 12'h777, 12'h666, 12'h777, 12'h777, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h988, 12'hDAA, 12'hC88, 12'hC88, 12'hD88, 12'hEAA, 12'hE99, 12'hD99, 12'hEAA, 12'hFBB, 12'hFBB, 12'hEBA, 12'hD99, 12'hC99, 12'hDA9, 12'hCA9, 12'hEBA, 12'hEBB, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hB87, 12'hB87, 12'hC88, 12'hB88, 12'hB88, 12'hA77, 12'h977, 12'h977, 12'h644, 12'h644, 12'h544, 12'h866, 12'h855, 12'hA76, 12'hA67, 12'h955, 12'h955, 12'hA55, 12'hB77, 12'hB66, 12'hC77, 12'hD99, 12'hD99, 12'hC98, 12'hD99, 12'hD99, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hC99, 12'hB88, 12'h966, 12'h744, 12'h633, 12'h532, 12'h422, 12'h422, 12'h533, 12'h533, 12'h644, 12'h644, 12'h644, 12'h644, 12'h745, 12'h533, 12'h756, 12'h755, 12'h645, 12'h211, 12'h433, 12'h533, 12'h534, 12'h533, 12'h423, 12'h422, 12'h533, 12'h533, 12'h533, 12'h633, 12'h533, 12'h533, 12'h533, 12'h543, 12'h544, 12'h544, 12'h533, 12'h533, 12'h433, 12'h433, 12'h544, 12'h544, 12'h333, 12'h433, 12'h655, 12'h655, 12'h555, 12'h766, 12'h878, 12'h777, 12'h878, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h667, 12'h776, 12'h677, 12'h767, 12'h676, 12'h767, 12'h776, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h777, 12'h778, 12'h777, 12'h777, 12'h776, 12'h866, 12'h977, 12'hC99, 12'hC88, 12'hC88, 12'hD99, 12'hEAA, 12'hE99, 12'hD99, 12'hEBB, 12'hFBB, 12'hFBB, 12'hFBA, 12'hEBA, 12'hC98, 12'hDA9, 12'hDA9, 12'hEAA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBA, 12'hDAA, 12'hEBA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hD9A, 12'hC99, 12'hD99, 12'hC99, 12'hB88, 12'hB77, 12'hA77, 12'h966, 12'h965, 12'h966, 12'hA66, 12'hA66, 12'hA66, 12'hB77, 12'hB77, 12'hC88, 12'hD99, 12'hDA9, 12'hDA9, 12'hDAA, 12'hD99, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hC98, 12'hB87, 12'h966, 12'h744, 12'h533, 12'h532, 12'h532, 12'h533, 12'h643, 12'h633, 12'h422, 12'h523, 12'h634, 12'h755, 12'h977, 12'h644, 12'h756, 12'h433, 12'h211, 12'h222, 12'h544, 12'h545, 12'h755, 12'h655, 12'h533, 12'h422, 12'h422, 12'h422, 12'h432, 12'h533, 12'h533, 12'h433, 12'h533, 12'h544, 12'h544, 12'h544, 12'h533, 12'h433, 12'h534, 12'h433, 12'h544, 12'h544, 12'h423, 12'h322, 12'h433, 12'h534, 12'h534, 12'h534, 12'h655, 12'h877, 12'h766, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h788,
		12'h666, 12'h666, 12'h666, 12'h676, 12'h777, 12'h677, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h877, 12'h977, 12'hDAA, 12'hD9A, 12'hE9A, 12'hE99, 12'hE99, 12'hFAA, 12'hEAA, 12'hEBA, 12'hEBA, 12'hFBA, 12'hEB9, 12'hDA9, 12'hDA9, 12'hDBA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hDBB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBA, 12'hEAA, 12'hDAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC98, 12'hC88, 12'hD99, 12'hC88, 12'hC88, 12'hC88, 12'hB77, 12'hB77, 12'hB77, 12'hB76, 12'hB66, 12'hB76, 12'hB77, 12'hB77, 12'hC88, 12'hC88, 12'hC98, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hEAA, 12'hEAA, 12'hD99, 12'hD88, 12'hB78, 12'hB77, 12'h855, 12'h744, 12'h643, 12'h533, 12'h533, 12'h633, 12'h644, 12'h634, 12'h744, 12'h844, 12'h855, 12'h855, 12'h966, 12'h967, 12'h967, 12'h966, 12'h855, 12'h755, 12'h745, 12'h744, 12'h744, 12'h644, 12'h644, 12'h633, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h533, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h433, 12'h433, 12'h433, 12'h534, 12'h544, 12'h433, 12'h422, 12'h533, 12'h422, 12'h311, 12'h211, 12'h544, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h677, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h787, 12'h888, 12'h777, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h866, 12'hB99, 12'hEBB, 12'hE9A, 12'hE99, 12'hE99, 12'hFBB, 12'hEA9, 12'hDA9, 12'hEA9, 12'hEA9, 12'hC98, 12'hA76, 12'hDA9, 12'hEBA, 12'hDA9, 12'hDAA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hECB, 12'hEBB, 12'hECB, 12'hECC, 12'hECB, 12'hEBB, 12'hEBB, 12'hECB, 12'hECB, 12'hEBB, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hEA9, 12'hDA9, 12'hEAA, 12'hDA9, 12'hD99, 12'hEAA, 12'hD99, 12'hD98, 12'hC98, 12'hC88, 12'hC88, 12'hC88, 12'hC77, 12'hC77, 12'hC77, 12'hC88, 12'hC88, 12'hC88, 12'hC98, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD9A, 12'hE99, 12'hEAA, 12'hE99, 12'hC88, 12'hC78, 12'hB77, 12'h855, 12'h744, 12'h634, 12'h533, 12'h644, 12'h644, 12'h633, 12'h644, 12'h744, 12'h744, 12'h845, 12'h845, 12'h955, 12'hA66, 12'hA77, 12'hA77, 12'hA76, 12'hA67, 12'h966, 12'h966, 12'h866, 12'h855, 12'h755, 12'h755, 12'h644, 12'h644, 12'h643, 12'h543, 12'h533, 12'h543, 12'h644, 12'h643, 12'h644, 12'h543, 12'h533, 12'h433, 12'h533, 12'h533, 12'h433, 12'h433, 12'h432, 12'h422, 12'h422, 12'h211, 12'h311, 12'h211, 12'h666, 12'h887, 12'h888, 12'h887, 12'h877, 12'h877, 12'h877, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h676, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h777, 12'h788, 12'h787, 12'h877, 12'h888, 12'h777, 12'h887, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h777, 12'h777, 12'h877, 12'h866, 12'hC99, 12'hDAA, 12'hE99, 12'hFAA, 12'hFBB, 12'hE99, 12'hD98, 12'hE99, 12'hE98, 12'hC98, 12'hB87, 12'hEBA, 12'hFCB, 12'hDA9, 12'hDAA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hECB, 12'hEBB, 12'hEBB, 12'hECB, 12'hEBB, 12'hEBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hEAA, 12'hEAA, 12'hD99, 12'hDA9, 12'hEAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC98, 12'hC88, 12'hC88, 12'hD98, 12'hD99, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD98, 12'hD89, 12'hD99, 12'hD99, 12'hD99, 12'hE99, 12'hD99, 12'hC88, 12'hC88, 12'hB77, 12'h854, 12'h644, 12'h634, 12'h633, 12'h644, 12'h744, 12'h744, 12'h634, 12'h744, 12'h855, 12'h744, 12'h744, 12'h844, 12'h845, 12'h844, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h744, 12'h744, 12'h744, 12'h644, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h654, 12'h644, 12'h644, 12'h544, 12'h533, 12'h433, 12'h434, 12'h433, 12'h422, 12'h433, 12'h422, 12'h322, 12'h422, 12'h311, 12'h322, 12'h433, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777,
		12'h667, 12'h776, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h788, 12'h778, 12'h887, 12'h788, 12'h777, 12'h878, 12'h788, 12'h777, 12'h878, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h877, 12'h977, 12'hDAA, 12'hEAA, 12'hFAB, 12'hFAA, 12'hE99, 12'hE99, 12'hD98, 12'hD99, 12'hD98, 12'hEBA, 12'hFDB, 12'hFCB, 12'hDA9, 12'hDA9, 12'hDBA, 12'hEBA, 12'hEBB, 12'hECB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hEBB, 12'hECB, 12'hECB, 12'hFCC, 12'hFCB, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEAA, 12'hDAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC88, 12'hC98, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hEAA, 12'hEAA, 12'hEA9, 12'hD99, 12'hD99, 12'hD99, 12'hD98, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hE9A, 12'hD99, 12'hD99, 12'hC88, 12'hB77, 12'h844, 12'h644, 12'h633, 12'h533, 12'h644, 12'h644, 12'h744, 12'h744, 12'h744, 12'h855, 12'h956, 12'h966, 12'h955, 12'h855, 12'h855, 12'h855, 12'h955, 12'h955, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h866, 12'h865, 12'h855, 12'h755, 12'h755, 12'h754, 12'h755, 12'h654, 12'h644, 12'h544, 12'h533, 12'h433, 12'h433, 12'h423, 12'h433, 12'h422, 12'h422, 12'h533, 12'h312, 12'h432, 12'h766, 12'h988, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h877, 12'h777, 12'h777, 12'h787, 12'h777, 12'h877, 12'h787, 12'h777, 12'h777,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h787, 12'h778, 12'h888, 12'h877, 12'h777, 12'h777, 12'h888, 12'h787, 12'h878, 12'h888, 12'h787, 12'h877, 12'h878, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h876, 12'hCAA, 12'hEBB, 12'hFBB, 12'hEAA, 12'hD88, 12'hD88, 12'hE99, 12'hEAA, 12'hEBA, 12'hFCB, 12'hFCB, 12'hECB, 12'hDBA, 12'hDAA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hECB, 12'hECB, 12'hDBB, 12'hDBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hECB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEAA, 12'hEAA, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hEAA, 12'hD99, 12'hEAA, 12'hE9A, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hD99, 12'hD99, 12'hD99, 12'hD9A, 12'hD99, 12'hD99, 12'hD99, 12'hC88, 12'hB77, 12'hA66, 12'h855, 12'h634, 12'h633, 12'h644, 12'h644, 12'h634, 12'h634, 12'h744, 12'h844, 12'h855, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h955, 12'h865, 12'h865, 12'h966, 12'h966, 12'h865, 12'h855, 12'h855, 12'h754, 12'h644, 12'h644, 12'h644, 12'h433, 12'h534, 12'h433, 12'h433, 12'h422, 12'h422, 12'h433, 12'h633, 12'h423, 12'h544, 12'h877, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h887, 12'h888,
		12'h676, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h778, 12'h777, 12'h787, 12'h878, 12'h787, 12'h777, 12'h778, 12'h787, 12'h877, 12'h788, 12'h888, 12'h777, 12'h787, 12'h778, 12'h777, 12'h777, 12'h777, 12'h877, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h876, 12'hB99, 12'hDAA, 12'hFBB, 12'hFAA, 12'hC78, 12'hD88, 12'hE99, 12'hFBA, 12'hEBA, 12'hDAA, 12'hEBB, 12'hECB, 12'hDBA, 12'hEAA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hECB, 12'hEBB, 12'hEBA, 12'hDBA, 12'hDBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hE9A, 12'hD99, 12'hD99, 12'hD99, 12'hE9A, 12'hD89, 12'hC88, 12'hB77, 12'hA66, 12'h855, 12'h633, 12'h633, 12'h634, 12'h644, 12'h633, 12'h644, 12'h744, 12'h744, 12'h845, 12'h855, 12'h955, 12'h956, 12'h956, 12'h956, 12'h966, 12'h956, 12'h956, 12'h956, 12'h966, 12'h956, 12'h966, 12'h966, 12'h966, 12'h966, 12'h966, 12'h966, 12'h865, 12'h966, 12'h966, 12'h865, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h533, 12'h423, 12'h433, 12'h422, 12'h422, 12'h533, 12'h543, 12'h533, 12'h655, 12'h877, 12'h888, 12'h787, 12'h888, 12'h888, 12'h887, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887,
		12'h777, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h778, 12'h877, 12'h777, 12'h787, 12'h788, 12'h777, 12'h788, 12'h888, 12'h877, 12'h788, 12'h888, 12'h878, 12'h777, 12'h787, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h777, 12'h777, 12'h777, 12'h877, 12'h877, 12'hA88, 12'hDAA, 12'hFBB, 12'hFBB, 12'hD99, 12'hB77, 12'hC78, 12'hE99, 12'hFBB, 12'hDAA, 12'hEBB, 12'hFCB, 12'hDAA, 12'hDBA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBB, 12'hDBA, 12'hDBA, 12'hEBA, 12'hEBB, 12'hECB, 12'hFBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hEAA, 12'hDAA, 12'hEAA, 12'hD9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hE99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hE99, 12'hD99, 12'hDAA, 12'hD99, 12'hD9A, 12'hD99, 12'hD99, 12'hE9A, 12'hD99, 12'hC88, 12'hB77, 12'hB77, 12'h855, 12'h744, 12'h644, 12'h643, 12'h634, 12'h644, 12'h734, 12'h744, 12'h744, 12'h845, 12'h845, 12'h855, 12'h955, 12'h966, 12'h966, 12'h966, 12'h966, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA76, 12'hA66, 12'h966, 12'h855, 12'h754, 12'h855, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h433, 12'h423, 12'h422, 12'h422, 12'h423, 12'h533, 12'h533, 12'h544, 12'h755, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h788, 12'h777, 12'h777, 12'h888, 12'h777, 12'h877, 12'h878, 12'h787, 12'h888, 12'h778, 12'h887, 12'h888, 12'h888, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h867, 12'h777, 12'h777, 12'h877, 12'h877, 12'h877, 12'h977, 12'hEBB, 12'hD9A, 12'hDAA, 12'hFBB, 12'hFCB, 12'hEAA, 12'hD89, 12'hC98, 12'hC99, 12'hDAA, 12'hECB, 12'hDAA, 12'hEAA, 12'hEBA, 12'hEBA, 12'hEBB, 12'hDBA, 12'hDBA, 12'hEBB, 12'hDBA, 12'hDBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hECB, 12'hFBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hD9A, 12'hD99, 12'hD99, 12'hD9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD9A, 12'hE99, 12'hE9A, 12'hE99, 12'hE99, 12'hE9A, 12'hE9A, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD9A, 12'hD99, 12'hE99, 12'hD99, 12'hC88, 12'hC77, 12'hB77, 12'h955, 12'h744, 12'h644, 12'h644, 12'h644, 12'h744, 12'h634, 12'h734, 12'h744, 12'h844, 12'h845, 12'h845, 12'h955, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h966, 12'h966, 12'h955, 12'h855, 12'h754, 12'h754, 12'h744, 12'h644, 12'h644, 12'h644, 12'h433, 12'h423, 12'h433, 12'h422, 12'h322, 12'h522, 12'h533, 12'h533, 12'h644, 12'h766, 12'h887, 12'h887, 12'h888, 12'h898, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h999, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h878, 12'h877, 12'h787, 12'h878, 12'h788, 12'h777, 12'h877, 12'h788, 12'h787, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h777, 12'h777, 12'h877, 12'h877, 12'h877, 12'h878, 12'h777, 12'h877, 12'h877, 12'h877, 12'hCAA, 12'hEBB, 12'hCAA, 12'hFCB, 12'hFBB, 12'hEBB, 12'hEAA, 12'hEAA, 12'hEBA, 12'hFBB, 12'hEBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hD99, 12'hD99, 12'hE9A, 12'hE9A, 12'hEAA, 12'hE99, 12'hD99, 12'hD9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hDAA, 12'hD9A, 12'hD9A, 12'hDAA, 12'hDAA, 12'hD99, 12'hC89, 12'hC88, 12'hB78, 12'h966, 12'h745, 12'h744, 12'h644, 12'h643, 12'h744, 12'h744, 12'h643, 12'h744, 12'h744, 12'h844, 12'h855, 12'h955, 12'h955, 12'h955, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hB66, 12'hB66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h855, 12'h755, 12'h755, 12'h744, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h432, 12'h422, 12'h422, 12'h523, 12'h533, 12'h633, 12'h644, 12'h534, 12'hA99, 12'h988, 12'h898, 12'h898, 12'h898, 12'h898, 12'h888, 12'h898, 12'h998, 12'h998, 12'h888, 12'h999, 12'h999, 12'h888, 12'h998, 12'h999, 12'h998, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h788, 12'h887, 12'h878, 12'h787, 12'h877, 12'h888, 12'h788, 12'h777, 12'h888, 12'h888, 12'h888, 12'h788, 12'h787, 12'h878, 12'h777, 12'h787, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h778, 12'h878, 12'h878, 12'h878, 12'h877, 12'h877, 12'hA88, 12'hDBB, 12'hECB, 12'hECB, 12'hEAA, 12'hDAA, 12'hDAA, 12'hEBB, 12'hEBA, 12'hEBA, 12'hEBA, 12'hDAA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBB, 12'hEBA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hD9A, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hC99, 12'hD99, 12'hD99, 12'hD9A, 12'hDAA, 12'hD99, 12'hDAA, 12'hDAA, 12'hEBB, 12'hDAA, 12'hD9A, 12'hC99, 12'hB78, 12'h966, 12'h855, 12'h744, 12'h744, 12'h634, 12'h633, 12'h633, 12'h633, 12'h744, 12'h744, 12'h744, 12'h854, 12'h855, 12'h955, 12'h955, 12'h956, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hB76, 12'hA67, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h965, 12'h855, 12'h755, 12'h744, 12'h744, 12'h644, 12'h544, 12'h644, 12'h544, 12'h543, 12'h433, 12'h433, 12'h433, 12'h533, 12'h533, 12'h634, 12'h644, 12'h655, 12'hA99, 12'h988, 12'h898, 12'h898, 12'h898, 12'h898, 12'h998, 12'h999, 12'h998, 12'h999, 12'h899, 12'h888, 12'h988, 12'h899, 12'h888, 12'h989, 12'h898, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h788, 12'h878, 12'h888, 12'h787, 12'h878, 12'h888, 12'h787, 12'h878, 12'h787, 12'h878, 12'h887, 12'h888, 12'h878, 12'h787, 12'h778, 12'h877, 12'h777, 12'h777, 12'h777, 12'h877, 12'h878, 12'h777, 12'h877, 12'h878, 12'h888, 12'h878, 12'h877, 12'h977, 12'hB99, 12'hFDD, 12'hFCC, 12'hFCC, 12'hEBA, 12'hDAA, 12'hEAA, 12'hEBA, 12'hEBB, 12'hEBB, 12'hEAA, 12'hDAA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hDBB, 12'hDBA, 12'hDBB, 12'hEBB, 12'hEBA, 12'hEBB, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAB, 12'hEBA, 12'hEBA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hD99, 12'hD99, 12'hD99, 12'hE99, 12'hD99, 12'hD99, 12'hD89, 12'hD88, 12'hC88, 12'hD88, 12'hC88, 12'hC88, 12'hD88, 12'hD89, 12'hC88, 12'hC88, 12'hD89, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hEBB, 12'hEBB, 12'hDAA, 12'hC89, 12'hB78, 12'hA66, 12'h855, 12'h744, 12'h744, 12'h644, 12'h633, 12'h633, 12'h633, 12'h644, 12'h744, 12'h744, 12'h844, 12'h855, 12'h955, 12'h955, 12'h955, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA76, 12'hA67, 12'hA66, 12'hA66, 12'h966, 12'h966, 12'h855, 12'h855, 12'h744, 12'h744, 12'h644, 12'h644, 12'h544, 12'h544, 12'h533, 12'h533, 12'h433, 12'h433, 12'h422, 12'h533, 12'h533, 12'h634, 12'h644, 12'h877, 12'h999, 12'h988, 12'h999, 12'h899, 12'h888, 12'h899, 12'h998, 12'h988, 12'h889, 12'h998, 12'h999, 12'h888, 12'h998, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h887, 12'h778, 12'h887, 12'h888, 12'h788, 12'h877, 12'h888, 12'h888, 12'h777, 12'h788, 12'h787, 12'h777, 12'h778, 12'h887, 12'h777, 12'h778, 12'h877, 12'h777, 12'h778, 12'h877, 12'h877, 12'h878, 12'h878, 12'h877, 12'h788, 12'h888, 12'h888, 12'h877, 12'h988, 12'h978, 12'hDCB, 12'hECC, 12'hFCC, 12'hFCC, 12'hFCB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hEBB, 12'hDBA, 12'hDAA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hEBB, 12'hEBA, 12'hDBB, 12'hEBB, 12'hEBA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hE9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC88, 12'hC78, 12'hB77, 12'hB77, 12'hB67, 12'hB67, 12'hB77, 12'hC77, 12'hC78, 12'hC88, 12'hD88, 12'hD89, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDAA, 12'hDAA, 12'hDAB, 12'hEAB, 12'hDAA, 12'hDAA, 12'hC89, 12'hB88, 12'hA66, 12'h845, 12'h845, 12'h744, 12'h644, 12'h644, 12'h634, 12'h633, 12'h633, 12'h633, 12'h634, 12'h744, 12'h845, 12'h855, 12'h855, 12'h955, 12'h965, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h956, 12'h855, 12'h744, 12'h744, 12'h755, 12'h644, 12'h644, 12'h633, 12'h544, 12'h543, 12'h533, 12'h433, 12'h422, 12'h422, 12'h533, 12'h633, 12'h633, 12'h644, 12'h988, 12'h988, 12'h988, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h988, 12'h888, 12'h898, 12'h988, 12'h889, 12'h898, 12'h988, 12'h888, 12'h998, 12'h989, 12'h888, 12'h888,
		12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h787, 12'h888, 12'h777, 12'h777, 12'h877, 12'h777, 12'h878, 12'h878, 12'h777, 12'h778, 12'h778, 12'h878, 12'h777, 12'h877, 12'h877, 12'hCBB, 12'hECC, 12'hFCC, 12'hFCC, 12'hFCC, 12'hFBB, 12'hEBB, 12'hDA9, 12'hDAA, 12'hDAA, 12'hEBA, 12'hEBA, 12'hEBA, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDAA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hEAA, 12'hEA9, 12'hD99, 12'hC88, 12'hC78, 12'hC77, 12'hA66, 12'hA66, 12'hA56, 12'hA66, 12'hB76, 12'hC77, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hD89, 12'hD99, 12'hE99, 12'hD99, 12'hD9A, 12'hDAA, 12'hE99, 12'hD9A, 12'hEAA, 12'hDAA, 12'hEAA, 12'hDAB, 12'hDAA, 12'hD99, 12'hC89, 12'hB77, 12'hA66, 12'h966, 12'h855, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h633, 12'h633, 12'h633, 12'h633, 12'h744, 12'h844, 12'h855, 12'h855, 12'h955, 12'h966, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h956, 12'h855, 12'h755, 12'h744, 12'h644, 12'h544, 12'h533, 12'h533, 12'h544, 12'h533, 12'h433, 12'h432, 12'h311, 12'h311, 12'h533, 12'h533, 12'h644, 12'h655, 12'h999, 12'h999, 12'h988, 12'h888, 12'h898, 12'h888, 12'h888, 12'h988, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h899, 12'h998, 12'h888, 12'h888,
		12'h888, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h788, 12'h877, 12'h777, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h887, 12'h788, 12'h878, 12'h887, 12'h877, 12'h877, 12'h887, 12'h888, 12'h878, 12'h788, 12'h778, 12'h888, 12'h877, 12'h878, 12'h877, 12'hDBB, 12'hDBB, 12'hEBB, 12'hEBB, 12'hDAA, 12'hD99, 12'hB87, 12'hC99, 12'hEAA, 12'hDBA, 12'hEBA, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hEAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hC88, 12'hC88, 12'hB88, 12'hB67, 12'hA66, 12'hA66, 12'hA66, 12'hB77, 12'hC77, 12'hC88, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hD89, 12'hD88, 12'hC88, 12'hB77, 12'hA66, 12'hB67, 12'hC88, 12'hD88, 12'hD99, 12'hEAA, 12'hD9A, 12'hEAA, 12'hEBB, 12'hEBB, 12'hDAA, 12'hC99, 12'hC88, 12'hB78, 12'hA67, 12'h855, 12'h754, 12'h644, 12'h633, 12'h533, 12'h533, 12'h533, 12'h522, 12'h422, 12'h633, 12'h633, 12'h533, 12'h623, 12'h633, 12'h744, 12'h844, 12'h845, 12'h955, 12'h956, 12'h966, 12'h966, 12'h966, 12'h966, 12'h956, 12'h855, 12'h855, 12'h744, 12'h644, 12'h644, 12'h533, 12'h533, 12'h543, 12'h544, 12'h533, 12'h433, 12'h422, 12'h422, 12'h433, 12'h533, 12'h544, 12'h644, 12'h755, 12'h999, 12'h998, 12'h888, 12'h898, 12'h898, 12'h888, 12'h988, 12'h988, 12'h988, 12'h988, 12'h898, 12'h898, 12'h999, 12'h999, 12'h988, 12'h898, 12'h889, 12'h888, 12'h888, 12'h888,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h777, 12'h888, 12'h777, 12'h888, 12'h878, 12'h777, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h878, 12'h887, 12'h878, 12'h788, 12'h888, 12'h878, 12'h877, 12'h888, 12'h887, 12'h878, 12'h788, 12'h888, 12'h878, 12'h888, 12'h878, 12'h878, 12'h978, 12'hA89, 12'hC99, 12'hC89, 12'hB88, 12'hA77, 12'h966, 12'hC99, 12'hDAA, 12'hDBA, 12'hDBB, 12'hEBB, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hEAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hEAA, 12'hEAA, 12'hDA9, 12'hD99, 12'hC99, 12'hB77, 12'hA66, 12'h955, 12'hA77, 12'hC88, 12'hC88, 12'hC88, 12'hC98, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hD89, 12'hD99, 12'hD89, 12'hD89, 12'hD99, 12'hD99, 12'hC88, 12'hC78, 12'hC88, 12'hD99, 12'hD88, 12'hD88, 12'hD89, 12'hD89, 12'hD9A, 12'hEAA, 12'hD99, 12'hC89, 12'hC88, 12'hC88, 12'hB78, 12'h856, 12'h644, 12'h633, 12'h433, 12'h311, 12'h311, 12'h311, 12'h311, 12'h412, 12'h422, 12'h533, 12'h633, 12'h633, 12'h633, 12'h633, 12'h633, 12'h623, 12'h733, 12'h744, 12'h855, 12'h955, 12'h955, 12'h956, 12'h956, 12'h855, 12'h855, 12'h755, 12'h744, 12'h634, 12'h533, 12'h533, 12'h433, 12'h433, 12'h533, 12'h533, 12'h422, 12'h322, 12'h422, 12'h533, 12'h533, 12'h533, 12'h533, 12'h877, 12'h999, 12'h888, 12'h898, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h888, 12'h998, 12'h999, 12'h988, 12'h888, 12'h888,
		12'h888, 12'h878, 12'h878, 12'h877, 12'h878, 12'h877, 12'h877, 12'h778, 12'h887, 12'h877, 12'h888, 12'h888, 12'h878, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h777, 12'h887, 12'h788, 12'h777, 12'h877, 12'h788, 12'h777, 12'h888, 12'h778, 12'h777, 12'h888, 12'h888, 12'h787, 12'h777, 12'h777, 12'h887, 12'h887, 12'h877, 12'h877, 12'h877, 12'h977, 12'h977, 12'h976, 12'h977, 12'hDAA, 12'hDBA, 12'hDAA, 12'hEAA, 12'hDBA, 12'hDBA, 12'hEBB, 12'hDBB, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDBA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hEAA, 12'hEAA, 12'hDA9, 12'hD99, 12'hD98, 12'hA76, 12'h965, 12'hA76, 12'hC99, 12'hC98, 12'hC88, 12'hC98, 12'hC88, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hD99, 12'hD89, 12'hC88, 12'hC78, 12'hC77, 12'hC88, 12'hC78, 12'hC77, 12'hC88, 12'hC88, 12'hD99, 12'hC89, 12'hB78, 12'hB78, 12'hB78, 12'h977, 12'h744, 12'h522, 12'h422, 12'h311, 12'h211, 12'h312, 12'h312, 12'h422, 12'h422, 12'h533, 12'h634, 12'h633, 12'h634, 12'h644, 12'h634, 12'h744, 12'h744, 12'h633, 12'h744, 12'h744, 12'h844, 12'h956, 12'h966, 12'h955, 12'h855, 12'h745, 12'h744, 12'h644, 12'h634, 12'h533, 12'h433, 12'h433, 12'h533, 12'h433, 12'h433, 12'h423, 12'h422, 12'h533, 12'h533, 12'h544, 12'h433, 12'h433, 12'h888, 12'h998, 12'h888, 12'h988, 12'h898, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h988, 12'h898, 12'h888, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h878, 12'h877, 12'h887, 12'h878, 12'h877, 12'h877, 12'h777, 12'h777, 12'h878, 12'h777, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h878, 12'h777, 12'h887, 12'h777, 12'h787, 12'h887, 12'h888, 12'h777, 12'h887, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h777, 12'h887, 12'h877, 12'h778, 12'h878, 12'h877, 12'h877, 12'h987, 12'hCBA, 12'hDBA, 12'hDAA, 12'hEBA, 12'hEBA, 12'hDBA, 12'hDBB, 12'hEBB, 12'hDBA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hC98, 12'hC88, 12'hA66, 12'hC98, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hE9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD88, 12'hD88, 12'hC88, 12'hC88, 12'hC78, 12'hB77, 12'hB77, 12'hA66, 12'hA67, 12'hA66, 12'h855, 12'h866, 12'h866, 12'h745, 12'h523, 12'h312, 12'h312, 12'h311, 12'h312, 12'h422, 12'h422, 12'h423, 12'h533, 12'h533, 12'h533, 12'h633, 12'h644, 12'h744, 12'h744, 12'h744, 12'h744, 12'h744, 12'h745, 12'h845, 12'h744, 12'h855, 12'h855, 12'h855, 12'h855, 12'h744, 12'h644, 12'h634, 12'h533, 12'h533, 12'h433, 12'h533, 12'h433, 12'h433, 12'h423, 12'h422, 12'h422, 12'h423, 12'h534, 12'h544, 12'h544, 12'h544, 12'h998, 12'h998, 12'h998, 12'h888, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h888, 12'h998, 12'h998, 12'h989, 12'h998, 12'h898, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h878, 12'h877, 12'h888, 12'h877, 12'h877, 12'h888, 12'h777, 12'h777, 12'h877, 12'h777, 12'h777, 12'h888, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h788, 12'h878, 12'h888, 12'h778, 12'h877, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h987, 12'hCBA, 12'hDA9, 12'hDA9, 12'hDBA, 12'hEAA, 12'hDBA, 12'hDBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hEAA, 12'hDBA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hC98, 12'hC87, 12'hB76, 12'hEA9, 12'hDA9, 12'hD99, 12'hDA9, 12'hC98, 12'hC99, 12'hDAA, 12'hDA9, 12'hDAA, 12'hD9A, 12'hE99, 12'hD9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC89, 12'hC78, 12'hB77, 12'hB77, 12'h955, 12'h844, 12'h844, 12'h744, 12'h744, 12'h633, 12'h633, 12'h533, 12'h522, 12'h422, 12'h422, 12'h523, 12'h533, 12'h533, 12'h533, 12'h534, 12'h634, 12'h634, 12'h634, 12'h644, 12'h644, 12'h644, 12'h744, 12'h745, 12'h755, 12'h855, 12'h855, 12'h855, 12'h744, 12'h744, 12'h865, 12'h855, 12'h755, 12'h644, 12'h533, 12'h433, 12'h422, 12'h433, 12'h434, 12'h433, 12'h433, 12'h322, 12'h312, 12'h533, 12'h433, 12'h534, 12'h544, 12'h533, 12'h655, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h898, 12'h888, 12'h998, 12'h988, 12'h898, 12'h998, 12'h999, 12'h899, 12'h989, 12'h999, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888,
		12'h877, 12'h878, 12'h877, 12'h877, 12'h778, 12'h877, 12'h777, 12'h777, 12'h877, 12'h877, 12'h778, 12'h887, 12'h778, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h777, 12'h887, 12'h777, 12'h787, 12'h888, 12'h777, 12'h778, 12'h888, 12'h777, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h987, 12'hCBA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hEBA, 12'hDBA, 12'hDBA, 12'hEBB, 12'hDBA, 12'hDAA, 12'hEBA, 12'hDA9, 12'hDAA, 12'hEB9, 12'hDA9, 12'hDA9, 12'hEA9, 12'hDA9, 12'hD98, 12'hC98, 12'hB87, 12'hEBA, 12'hEAA, 12'hDA9, 12'hD99, 12'hD99, 12'hC99, 12'hDA9, 12'hD99, 12'hDA9, 12'hDAA, 12'hE9A, 12'hDA9, 12'hD9A, 12'hE9A, 12'hD9A, 12'hD9A, 12'hE9A, 12'hD99, 12'hE9A, 12'hD99, 12'hD89, 12'hD89, 12'hC88, 12'hC78, 12'hB77, 12'hB67, 12'hA66, 12'h966, 12'h955, 12'h955, 12'h955, 12'h855, 12'h855, 12'h744, 12'h644, 12'h634, 12'h644, 12'h744, 12'h634, 12'h634, 12'h634, 12'h634, 12'h644, 12'h634, 12'h644, 12'h744, 12'h644, 12'h644, 12'h744, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h854, 12'h844, 12'h855, 12'h865, 12'h755, 12'h744, 12'h533, 12'h433, 12'h433, 12'h533, 12'h433, 12'h544, 12'h444, 12'h221, 12'h322, 12'h433, 12'h533, 12'h544, 12'h533, 12'h433, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h888, 12'h998, 12'h998, 12'h888, 12'h999, 12'h998, 12'h999, 12'h999, 12'h888, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888,
		12'h878, 12'h877, 12'h878, 12'h877, 12'h877, 12'h878, 12'h777, 12'h777, 12'h878, 12'h777, 12'h887, 12'h878, 12'h777, 12'h888, 12'h888, 12'h887, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h888, 12'h887, 12'h788, 12'h887, 12'h887, 12'h888, 12'h778, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h987, 12'hCBA, 12'hDBA, 12'hDA9, 12'hDA9, 12'hEBA, 12'hEBA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hEBA, 12'hDBA, 12'hDA9, 12'hEAA, 12'hDA9, 12'hDA9, 12'hEBA, 12'hDA9, 12'hD99, 12'hC98, 12'hC98, 12'hDA9, 12'hD98, 12'hD98, 12'hC98, 12'hC88, 12'hC88, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hEAA, 12'hEAA, 12'hE99, 12'hD99, 12'hEAA, 12'hE9A, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC88, 12'hC77, 12'hB67, 12'hB77, 12'hB77, 12'hC78, 12'hB67, 12'hA66, 12'hA66, 12'hA67, 12'hA67, 12'h956, 12'h955, 12'h845, 12'h845, 12'h744, 12'h745, 12'h745, 12'h744, 12'h744, 12'h644, 12'h644, 12'h744, 12'h744, 12'h744, 12'h855, 12'h966, 12'h956, 12'h956, 12'h855, 12'h855, 12'h844, 12'h744, 12'h855, 12'h966, 12'h966, 12'h755, 12'h533, 12'h422, 12'h433, 12'h534, 12'h433, 12'h332, 12'h433, 12'h666, 12'h322, 12'h322, 12'h222, 12'h433, 12'h655, 12'h888, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h889, 12'h898, 12'h888, 12'h888, 12'h888,
		12'h888, 12'h888, 12'h877, 12'h888, 12'h878, 12'h877, 12'h877, 12'h878, 12'h777, 12'h887, 12'h878, 12'h888, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h987, 12'hBA9, 12'hDBA, 12'hDA9, 12'hDA9, 12'hDAA, 12'hEBA, 12'hDBA, 12'hDBB, 12'hEAA, 12'hEBA, 12'hDAA, 12'hEBA, 12'hDB9, 12'hDAA, 12'hDAA, 12'hDB9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hC98, 12'hDA8, 12'hDA9, 12'hD99, 12'hC98, 12'hC88, 12'hC87, 12'hB87, 12'hB87, 12'hB87, 12'hB88, 12'hC88, 12'hC99, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD9A, 12'hD99, 12'hD89, 12'hD89, 12'hD99, 12'hD89, 12'hD88, 12'hC78, 12'hC88, 12'hC78, 12'hC77, 12'hB67, 12'hB77, 12'hB77, 12'hB77, 12'hB67, 12'hB67, 12'hA66, 12'h955, 12'h855, 12'h845, 12'h744, 12'h744, 12'h745, 12'h644, 12'h644, 12'h634, 12'h633, 12'h634, 12'h633, 12'h634, 12'h855, 12'h855, 12'h966, 12'h966, 12'h955, 12'h844, 12'h744, 12'h744, 12'h865, 12'hA77, 12'h966, 12'h755, 12'h422, 12'h433, 12'h533, 12'h544, 12'h433, 12'h333, 12'h544, 12'h999, 12'h999, 12'h888, 12'h888, 12'h988, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h899, 12'h998, 12'h889, 12'h999, 12'h999, 12'h998, 12'h989, 12'h999, 12'h998, 12'h888, 12'h898,
		12'h877, 12'h878, 12'h877, 12'h878, 12'h888, 12'h777, 12'h887, 12'h778, 12'h877, 12'h877, 12'h788, 12'h887, 12'h877, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h887, 12'hBA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDAA, 12'hEAA, 12'hDBA, 12'hDBA, 12'hEAA, 12'hEBA, 12'hDA9, 12'hEAA, 12'hEBA, 12'hEA9, 12'hEBA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD98, 12'hC98, 12'hC88, 12'hC88, 12'hB77, 12'h844, 12'h633, 12'h622, 12'h633, 12'h966, 12'hB87, 12'hA77, 12'h967, 12'hB77, 12'hA77, 12'hA66, 12'hA77, 12'hA77, 12'hA77, 12'hA67, 12'hA66, 12'hA77, 12'hA66, 12'hB77, 12'hB77, 12'hC78, 12'hB77, 12'hA67, 12'hA66, 12'h956, 12'h956, 12'h955, 12'h854, 12'h744, 12'h744, 12'h744, 12'h634, 12'h634, 12'h634, 12'h633, 12'h533, 12'h533, 12'h533, 12'h533, 12'h532, 12'h522, 12'h634, 12'h955, 12'h966, 12'h966, 12'h966, 12'h744, 12'h633, 12'h844, 12'hA76, 12'hA87, 12'h866, 12'h644, 12'h422, 12'h433, 12'h544, 12'h533, 12'h433, 12'h322, 12'h777, 12'h998, 12'h998, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h999, 12'h998, 12'h998, 12'h889, 12'h999, 12'h898, 12'h998, 12'h989, 12'h899, 12'h998, 12'h988,
		12'h878, 12'h877, 12'h887, 12'h877, 12'h878, 12'h877, 12'h888, 12'h777, 12'h878, 12'h888, 12'h778, 12'h878, 12'h888, 12'h788, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h888, 12'h888, 12'h987, 12'hBA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hEAA, 12'hDBA, 12'hDBA, 12'hEAA, 12'hEBA, 12'hDAA, 12'hDAA, 12'hEB9, 12'hDA9, 12'hEBA, 12'hEBA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD98, 12'hD98, 12'hC88, 12'hC88, 12'hC88, 12'hA77, 12'h955, 12'h733, 12'h633, 12'h866, 12'hECB, 12'hEBB, 12'hDBA, 12'hFDC, 12'hECC, 12'hCA9, 12'hDAA, 12'hFCC, 12'hDBA, 12'hB98, 12'hB99, 12'hCAA, 12'hB88, 12'hB77, 12'hA77, 12'h966, 12'h966, 12'h845, 12'h855, 12'h744, 12'h744, 12'h744, 12'h754, 12'h744, 12'h633, 12'h532, 12'h633, 12'h533, 12'h422, 12'h422, 12'h311, 12'h311, 12'h321, 12'h311, 12'h522, 12'h744, 12'h855, 12'h966, 12'hA66, 12'hA66, 12'h955, 12'h744, 12'h854, 12'h966, 12'hA76, 12'h976, 12'h644, 12'h532, 12'h432, 12'h544, 12'h544, 12'h533, 12'h433, 12'h333, 12'h998, 12'h999, 12'h888, 12'h999, 12'h998, 12'h988, 12'h999, 12'h999, 12'h9A9, 12'h9A9, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h988, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998,
		12'h888, 12'h887, 12'h878, 12'h788, 12'h877, 12'h887, 12'h778, 12'h887, 12'h887, 12'h887, 12'h877, 12'h888, 12'h787, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h987, 12'hA99, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDBA, 12'hDBA, 12'hDAA, 12'hDBA, 12'hEBA, 12'hDBA, 12'hDAA, 12'hDBA, 12'hEBA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hC98, 12'hC98, 12'hC88, 12'hC88, 12'hB87, 12'hC88, 12'hC88, 12'h966, 12'h744, 12'hB99, 12'hCBA, 12'hCA9, 12'hDBB, 12'hDBB, 12'hCBA, 12'hECB, 12'hFDD, 12'hECC, 12'hCBA, 12'hEDC, 12'hEDC, 12'hDCB, 12'hDBB, 12'hCA9, 12'h977, 12'hECC, 12'hDBA, 12'hBA9, 12'hB99, 12'h876, 12'hA87, 12'hBA9, 12'h987, 12'h755, 12'h755, 12'h755, 12'h543, 12'h433, 12'h422, 12'h200, 12'h200, 12'h210, 12'h422, 12'h755, 12'h866, 12'h966, 12'hA67, 12'hA77, 12'hA66, 12'h955, 12'h955, 12'hA77, 12'hB87, 12'h977, 12'h755, 12'h533, 12'h422, 12'h533, 12'h544, 12'h544, 12'h433, 12'h433, 12'h655, 12'hA99, 12'h998, 12'h9AA, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'hAA9, 12'hAA9, 12'h999, 12'hAA9, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h989, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999,
		12'h777, 12'h887, 12'h778, 12'h787, 12'h887, 12'h778, 12'h888, 12'h888, 12'h788, 12'h888, 12'h887, 12'h777, 12'h888, 12'h888, 12'h877, 12'h788, 12'h888, 12'h877, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h988, 12'h988, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDBA, 12'hEAA, 12'hDBA, 12'hEBA, 12'hDAA, 12'hDBA, 12'hEAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hC99, 12'hD99, 12'hD99, 12'hC99, 12'hC88, 12'hC88, 12'hD99, 12'hD99, 12'hD99, 12'hC88, 12'hA77, 12'h966, 12'h855, 12'hC98, 12'hB88, 12'h965, 12'hA77, 12'hCAA, 12'hCA9, 12'hCA9, 12'hECB, 12'hDCB, 12'hDDC, 12'hDBB, 12'hBA9, 12'hCAA, 12'hFDD, 12'hDCB, 12'hDBA, 12'hBA9, 12'hA88, 12'hCBB, 12'hBA9, 12'h876, 12'h866, 12'h766, 12'h644, 12'h533, 12'h533, 12'h422, 12'h311, 12'h532, 12'h744, 12'h855, 12'h966, 12'hA66, 12'hA66, 12'hA76, 12'hA66, 12'hA66, 12'hA66, 12'hA76, 12'hA77, 12'hA77, 12'h966, 12'h533, 12'h422, 12'h433, 12'h543, 12'h544, 12'h543, 12'h433, 12'h323, 12'h888, 12'hA99, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAA9, 12'hA99, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h898, 12'h999, 12'h998, 12'h999, 12'h998, 12'h998,
		12'h888, 12'h888, 12'h887, 12'h878, 12'h888, 12'h887, 12'h887, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h878, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h787, 12'h888, 12'h888, 12'h887, 12'h887, 12'h987, 12'hCAA, 12'hDA9, 12'hD99, 12'hD99, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDAA, 12'hEB9, 12'hDAA, 12'hDB9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hC99, 12'hD99, 12'hD99, 12'hD89, 12'hD89, 12'hC88, 12'hC78, 12'hB78, 12'hB77, 12'hB77, 12'hA66, 12'hB77, 12'hB77, 12'hB88, 12'hD99, 12'hC99, 12'hCA9, 12'hDAA, 12'hB88, 12'hDA9, 12'hEBB, 12'hDBA, 12'hC99, 12'hC99, 12'h855, 12'hA77, 12'h976, 12'h643, 12'h522, 12'h744, 12'h533, 12'h522, 12'h644, 12'h744, 12'h855, 12'h855, 12'h855, 12'h955, 12'hA66, 12'hA67, 12'hB67, 12'hA66, 12'hA66, 12'hA76, 12'hA76, 12'hA77, 12'hA77, 12'h966, 12'h744, 12'h422, 12'h422, 12'h533, 12'h544, 12'h543, 12'h433, 12'h322, 12'h444, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAA9, 12'hAA9, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998,
		12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h787, 12'h888, 12'h888, 12'h887, 12'h788, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h887, 12'h988, 12'hCAA, 12'hDA9, 12'hC99, 12'hC99, 12'hC99, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDBA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hEAA, 12'hD99, 12'hEAA, 12'hE9A, 12'hD89, 12'hD89, 12'hD89, 12'hD88, 12'hC78, 12'hC78, 12'hD89, 12'hC78, 12'hB77, 12'hC78, 12'hB67, 12'hB67, 12'hA66, 12'hB77, 12'hB67, 12'hB77, 12'hB67, 12'hA66, 12'hA66, 12'h955, 12'hA56, 12'h955, 12'h955, 12'h855, 12'h845, 12'h844, 12'h845, 12'h844, 12'h845, 12'h955, 12'hA66, 12'hA67, 12'hA66, 12'hA66, 12'hA76, 12'hA66, 12'hA77, 12'hA87, 12'h976, 12'h865, 12'h754, 12'h533, 12'h533, 12'h543, 12'h644, 12'h533, 12'h433, 12'h433, 12'h322, 12'h877, 12'hA99, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'hAA9, 12'hAA9, 12'h999, 12'h9A9, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h899, 12'h998, 12'h998, 12'h999, 12'h998, 12'h999, 12'h998, 12'h998,
		12'h887, 12'h878, 12'h788, 12'h887, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h988, 12'hDBB, 12'hCAA, 12'hDAA, 12'hDA9, 12'hC99, 12'hB98, 12'hB98, 12'hC99, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hE9A, 12'hDA9, 12'hD9A, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAA, 12'hEAB, 12'hEAA, 12'hE9A, 12'hD9A, 12'hD9A, 12'hD99, 12'hD89, 12'hD89, 12'hD89, 12'hC67, 12'hC77, 12'hB77, 12'hC78, 12'hB77, 12'hC77, 12'hA66, 12'hA66, 12'hA66, 12'h955, 12'h945, 12'h844, 12'h844, 12'h744, 12'h744, 12'h744, 12'h744, 12'h844, 12'h855, 12'h956, 12'h966, 12'h966, 12'h955, 12'h965, 12'hA66, 12'hA77, 12'h976, 12'h976, 12'h855, 12'h644, 12'h532, 12'h422, 12'h533, 12'h544, 12'h544, 12'h433, 12'h433, 12'h322, 12'h555, 12'h999, 12'h999, 12'hAAA, 12'hAA9, 12'hAA9, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h887, 12'h878, 12'h888, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h888, 12'h998, 12'h988, 12'hCBA, 12'hCAA, 12'hC99, 12'hCA9, 12'hC99, 12'hC98, 12'hB87, 12'hC98, 12'hC99, 12'hCA9, 12'hCA9, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hD99, 12'hDAA, 12'hDA9, 12'hE99, 12'hDA9, 12'hD99, 12'hD9A, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hD89, 12'hC88, 12'hC78, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hC78, 12'hB77, 12'hA67, 12'hA66, 12'hA66, 12'hA56, 12'h955, 12'h845, 12'h844, 12'h744, 12'h744, 12'h744, 12'h744, 12'h744, 12'h965, 12'h865, 12'h855, 12'h855, 12'h855, 12'h855, 12'h865, 12'h976, 12'h976, 12'h866, 12'h755, 12'h643, 12'h543, 12'h533, 12'h533, 12'h654, 12'h543, 12'h433, 12'h434, 12'h322, 12'h433, 12'h999, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAA9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h998, 12'h999, 12'h999, 12'h998, 12'h898, 12'h999, 12'h999, 12'h898, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h988, 12'h898, 12'h988, 12'h888, 12'h998, 12'h898, 12'h998, 12'h988, 12'hCBA, 12'hDBA, 12'hC99, 12'hCA9, 12'hC99, 12'hC98, 12'hC98, 12'hB98, 12'hB98, 12'hC98, 12'hC98, 12'hC98, 12'hC99, 12'hCA9, 12'hC99, 12'hD99, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hDA9, 12'hD9A, 12'hD99, 12'hDA9, 12'hD99, 12'hD9A, 12'hDAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hC88, 12'hC78, 12'hC78, 12'hB77, 12'hB77, 12'hB77, 12'hB78, 12'hB67, 12'hA66, 12'hA67, 12'hA67, 12'hA66, 12'h956, 12'h955, 12'h844, 12'h744, 12'h744, 12'h744, 12'h744, 12'h855, 12'h955, 12'h866, 12'h855, 12'h854, 12'h754, 12'h754, 12'h865, 12'h865, 12'h865, 12'h754, 12'h643, 12'h543, 12'h532, 12'h433, 12'h543, 12'h433, 12'h433, 12'h433, 12'h332, 12'h545, 12'h999, 12'h999, 12'h9A9, 12'hAAA, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h898, 12'h988, 12'h998, 12'h999, 12'h998, 12'h998, 12'h999,
		12'h888, 12'h777, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h898, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h888, 12'h998, 12'h888, 12'h999, 12'h998, 12'hCAA, 12'hDBB, 12'hCA9, 12'hDA9, 12'hC98, 12'hDA9, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB98, 12'hC98, 12'hC98, 12'hC98, 12'hCA9, 12'hCA9, 12'hD99, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hDA9, 12'hDA9, 12'hD99, 12'hEA9, 12'hD99, 12'hE99, 12'hEAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD88, 12'hC88, 12'hC78, 12'hC78, 12'hC88, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hA76, 12'h966, 12'h955, 12'h855, 12'h844, 12'h844, 12'h845, 12'h855, 12'h855, 12'h855, 12'h855, 12'h855, 12'h744, 12'h744, 12'h754, 12'h754, 12'h754, 12'h654, 12'h644, 12'h643, 12'h543, 12'h533, 12'h533, 12'h443, 12'h433, 12'h433, 12'h322, 12'h433, 12'hA99, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h9A9, 12'h9A9, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h998, 12'h998, 12'h999, 12'h998, 12'h998, 12'h999, 12'h998, 12'h998, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h898, 12'h998, 12'h889, 12'h898, 12'h998, 12'h989, 12'h998, 12'h998,
		12'h777, 12'h777, 12'h778, 12'h888, 12'h788, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h988, 12'h898, 12'h998, 12'h898, 12'h898, 12'h898, 12'h988, 12'h998, 12'h988, 12'hBAA, 12'hECC, 12'hDAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hC98, 12'hB88, 12'hB88, 12'hB87, 12'hB88, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hCA9, 12'hC99, 12'hCA9, 12'hDA9, 12'hDAA, 12'hDAA, 12'hEAA, 12'hDAA, 12'hEA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hDAA, 12'hE99, 12'hEAA, 12'hD99, 12'hD99, 12'hD99, 12'hD89, 12'hC88, 12'hC77, 12'hB77, 12'hB77, 12'hC77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hA77, 12'hA66, 12'hA66, 12'h955, 12'h955, 12'h956, 12'h955, 12'h854, 12'h955, 12'h855, 12'h844, 12'h855, 12'h854, 12'h754, 12'h744, 12'h755, 12'h865, 12'h744, 12'h644, 12'h544, 12'h544, 12'h533, 12'h433, 12'h433, 12'h543, 12'h433, 12'h332, 12'h222, 12'h332, 12'h998, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'hA99, 12'hAAA, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h998, 12'h999, 12'h998, 12'h998, 12'h998, 12'h998, 12'h998, 12'h998, 12'h999, 12'h998, 12'h989, 12'h999, 12'h889, 12'h898, 12'h999, 12'h988, 12'h998,
		12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h777, 12'h887, 12'h888, 12'h878, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h988, 12'h888, 12'h898, 12'h888, 12'h898, 12'h998, 12'h988, 12'h998, 12'h988, 12'hA99, 12'hDCB, 12'hDBB, 12'hDBA, 12'hC99, 12'hC99, 12'hDA9, 12'hC99, 12'hC98, 12'hC88, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB88, 12'hC98, 12'hC98, 12'hCA8, 12'hCA9, 12'hCA9, 12'hC99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hD98, 12'hC88, 12'hC88, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hB77, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h955, 12'h955, 12'h955, 12'h844, 12'h754, 12'h744, 12'h744, 12'h754, 12'h755, 12'h755, 12'h644, 12'h643, 12'h533, 12'h533, 12'h433, 12'h432, 12'h443, 12'h544, 12'h332, 12'h211, 12'h433, 12'h988, 12'hAAA, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h999, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h899, 12'h899, 12'h998, 12'h899, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h898, 12'h898, 12'h989, 12'h998, 12'h988, 12'h899, 12'h998, 12'h999,
		12'h878, 12'h788, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h778, 12'h888, 12'h887, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h988, 12'h888, 12'h999, 12'h889, 12'h998, 12'h989, 12'h888, 12'h898, 12'h888, 12'h989, 12'h998, 12'h988, 12'h999, 12'hDBB, 12'hDBB, 12'hEBB, 12'hC99, 12'hC98, 12'hC98, 12'hC99, 12'hC99, 12'hC98, 12'hC98, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB97, 12'hB98, 12'hC98, 12'hC98, 12'hC99, 12'hC99, 12'hC98, 12'hC99, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDAA, 12'hEAA, 12'hDA9, 12'hDAA, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hC99, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC77, 12'hB77, 12'hB77, 12'hB77, 12'hB66, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'hA66, 12'hA66, 12'hA66, 12'h966, 12'h966, 12'h965, 12'h855, 12'h744, 12'h744, 12'h744, 12'h755, 12'h755, 12'h644, 12'h533, 12'h533, 12'h433, 12'h433, 12'h543, 12'h433, 12'h433, 12'h322, 12'h222, 12'h766, 12'h999, 12'h9A9, 12'hAAA, 12'hAA9, 12'h999, 12'hAA9, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h898, 12'h999, 12'h998, 12'h898, 12'h998, 12'h988, 12'h898, 12'h898, 12'h998, 12'h899, 12'h898, 12'h999, 12'h988, 12'h899, 12'h998, 12'h989, 12'h899, 12'h998, 12'h988, 12'h999,
		12'h787, 12'h878, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h788, 12'h888, 12'h787, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h988, 12'h898, 12'h998, 12'h989, 12'h898, 12'h998, 12'h999, 12'h888, 12'h888, 12'h898, 12'h899, 12'h888, 12'h988, 12'hBAA, 12'hECC, 12'hDBB, 12'hDBB, 12'hDAA, 12'hDA9, 12'hD99, 12'hC99, 12'hDA9, 12'hC99, 12'hC98, 12'hC98, 12'hB87, 12'hB88, 12'hB87, 12'hB87, 12'hB88, 12'hB98, 12'hB98, 12'hC98, 12'hC98, 12'hC98, 12'hCA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hC99, 12'hD99, 12'hD89, 12'hC99, 12'hD98, 12'hD89, 12'hC88, 12'hC88, 12'hD89, 12'hC88, 12'hC77, 12'hC78, 12'hB77, 12'hB77, 12'hA66, 12'hA66, 12'hA66, 12'h965, 12'h966, 12'hA66, 12'hA66, 12'h966, 12'hA66, 12'h966, 12'h855, 12'h855, 12'h744, 12'h755, 12'h855, 12'h644, 12'h644, 12'h533, 12'h433, 12'h433, 12'h433, 12'h432, 12'h433, 12'h322, 12'h211, 12'h666, 12'hAAA, 12'h999, 12'h999, 12'h999, 12'h9AA, 12'hAA9, 12'hA9A, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h898, 12'h998, 12'h989, 12'h898, 12'h988, 12'h999, 12'h888, 12'h998, 12'h989, 12'h898, 12'h998, 12'h998, 12'h989, 12'h899, 12'h998, 12'h988, 12'h899, 12'h998, 12'h989, 12'h999,
		12'h888, 12'h777, 12'h887, 12'h778, 12'h777, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h998, 12'h998, 12'h999, 12'h999, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h999, 12'h999, 12'h898, 12'h889, 12'h888, 12'hDED, 12'hFEE, 12'hDBB, 12'hECB, 12'hDAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hDA9, 12'hCA9, 12'hC98, 12'hC98, 12'hC98, 12'hB98, 12'hB98, 12'hB88, 12'hB87, 12'hB87, 12'hB87, 12'hB98, 12'hB98, 12'hB98, 12'hB98, 12'hB99, 12'hC99, 12'hCA9, 12'hDAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hD99, 12'hC99, 12'hC99, 12'hD98, 12'hD99, 12'hD99, 12'hC88, 12'hC98, 12'hC98, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hB88, 12'hB88, 12'hB77, 12'hB77, 12'hA66, 12'hA66, 12'h965, 12'h955, 12'h966, 12'h955, 12'h855, 12'h844, 12'h744, 12'h744, 12'h744, 12'h744, 12'h644, 12'h643, 12'h533, 12'h533, 12'h433, 12'h432, 12'h433, 12'h332, 12'h222, 12'h433, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h898, 12'h999, 12'h999, 12'h898, 12'h989, 12'h998, 12'h899, 12'h988, 12'h999, 12'h998, 12'h889, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h878, 12'h787, 12'h888, 12'h888, 12'h878, 12'h888, 12'h878, 12'h888, 12'h878, 12'h888, 12'h878, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h898, 12'h988, 12'h898, 12'h888, 12'h989, 12'h899, 12'h998, 12'h989, 12'h988, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h988, 12'h999, 12'h999, 12'h999, 12'h898, 12'hAAA, 12'hFFF, 12'hFFE, 12'hEDD, 12'hCAA, 12'hDBA, 12'hDA9, 12'hC99, 12'hC98, 12'hDA9, 12'hDA9, 12'hD99, 12'hC98, 12'hC98, 12'hC98, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hA88, 12'hA88, 12'hB88, 12'hB98, 12'hC99, 12'hC99, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hEAA, 12'hEAA, 12'hDAA, 12'hD99, 12'hD99, 12'hDA9, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hC88, 12'hB77, 12'hB77, 12'hC88, 12'hC88, 12'hC88, 12'hB77, 12'hB77, 12'hB77, 12'hA77, 12'hA66, 12'hA66, 12'h955, 12'h965, 12'h855, 12'h855, 12'h744, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h533, 12'h433, 12'h432, 12'h322, 12'h322, 12'h332, 12'h333, 12'h777, 12'hAA9, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h889, 12'h898, 12'h989, 12'h998, 12'h898, 12'h989, 12'h998, 12'h898, 12'h988, 12'h899, 12'h998, 12'h989, 12'h899, 12'h998, 12'h999, 12'h988, 12'h998, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h777, 12'h888, 12'h888, 12'h787, 12'h878, 12'h787, 12'h887, 12'h788, 12'h777, 12'h888, 12'h777, 12'h788, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h998, 12'h899, 12'h989, 12'h998, 12'h899, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAAA, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hECC, 12'hDBB, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hC99, 12'hC99, 12'hC98, 12'hB98, 12'hB88, 12'hB98, 12'hA88, 12'hA88, 12'hA87, 12'hA88, 12'hB88, 12'hB98, 12'hB98, 12'hC99, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hEBA, 12'hEBA, 12'hEAA, 12'hDAA, 12'hDA9, 12'hD99, 12'hC99, 12'hC99, 12'hC88, 12'hC88, 12'hC88, 12'hB77, 12'hB77, 12'hC88, 12'hC88, 12'hC88, 12'hB77, 12'hB87, 12'hB77, 12'hA77, 12'hA66, 12'h966, 12'h966, 12'h855, 12'h755, 12'h744, 12'h644, 12'h644, 12'h644, 12'h644, 12'h543, 12'h433, 12'h432, 12'h322, 12'h322, 12'h322, 12'h333, 12'h121, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h989, 12'h898, 12'h998, 12'h889, 12'h998, 12'h999, 12'h998, 12'h998, 12'h999, 12'h998, 12'h999, 12'h999, 12'h899, 12'h999, 12'h998, 12'h989, 12'h999, 12'h999, 12'h999,
		12'h787, 12'h878, 12'h877, 12'h788, 12'h888, 12'h887, 12'h778, 12'h888, 12'h888, 12'h887, 12'h888, 12'h788, 12'h877, 12'h777, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h998, 12'h988, 12'h999, 12'h999, 12'h898, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hECB, 12'hDAA, 12'hDAA, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hCA9, 12'hC98, 12'hB98, 12'hB98, 12'hB88, 12'hB88, 12'hA87, 12'hA87, 12'hA87, 12'hA87, 12'hA88, 12'hB88, 12'hB98, 12'hC99, 12'hCA9, 12'hCA9, 12'hDA9, 12'hDAA, 12'hDA9, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hD99, 12'hD99, 12'hC99, 12'hC89, 12'hC88, 12'hB77, 12'hB88, 12'hC88, 12'hC88, 12'hC88, 12'hB88, 12'hC88, 12'hC88, 12'hB88, 12'hB88, 12'hB77, 12'hA66, 12'h966, 12'h966, 12'h855, 12'h754, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h332, 12'h221, 12'h898, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h989, 12'h898, 12'h998, 12'h999, 12'h998, 12'h999, 12'h888, 12'h998, 12'h899, 12'h989, 12'h898, 12'h999, 12'h998, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h878, 12'h888, 12'h778, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h999, 12'h999, 12'h889, 12'h898, 12'h998, 12'h988, 12'h888, 12'h999, 12'h999, 12'h998, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h777, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEDC, 12'hCBB, 12'hCA9, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hCA9, 12'hDA9, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hC98, 12'hB88, 12'hB98, 12'hB98, 12'hB88, 12'hA88, 12'hA88, 12'hB88, 12'hA88, 12'hA88, 12'hB98, 12'hB98, 12'hB99, 12'hC99, 12'hDA9, 12'hC99, 12'hC99, 12'hD99, 12'hD99, 12'hD99, 12'hC99, 12'hC98, 12'hC88, 12'hC88, 12'hC87, 12'hB77, 12'hB77, 12'hB77, 12'hB87, 12'hB77, 12'hB87, 12'hC88, 12'hB88, 12'hB88, 12'hA77, 12'hA76, 12'h966, 12'h966, 12'h855, 12'h755, 12'h644, 12'h533, 12'h533, 12'h544, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h332, 12'h767, 12'h999, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h899, 12'h888, 12'h999, 12'h899, 12'h989, 12'h999, 12'h898, 12'h999, 12'h999, 12'h999, 12'h899, 12'h999, 12'h999, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h888, 12'h787, 12'h888, 12'h888, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h988, 12'h999, 12'h999, 12'h989, 12'h899, 12'h999, 12'h998, 12'h998, 12'h999, 12'h998, 12'h898, 12'h999, 12'h999, 12'h999, 12'h888, 12'h666, 12'h9AA, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEDC, 12'hCAA, 12'hCAA, 12'hCAA, 12'hCA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD99, 12'hD98, 12'hC98, 12'hC98, 12'hB88, 12'hB88, 12'hB88, 12'hB98, 12'hB98, 12'hB98, 12'hA88, 12'hA87, 12'hA87, 12'hA87, 12'hA88, 12'hA88, 12'hB88, 12'hB98, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB98, 12'hB88, 12'hB88, 12'hB88, 12'hB88, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA77, 12'hA88, 12'hA77, 12'hA77, 12'h976, 12'h855, 12'h755, 12'h654, 12'h644, 12'h533, 12'h533, 12'h533, 12'h433, 12'h332, 12'h322, 12'h322, 12'h322, 12'h332, 12'h222, 12'h332, 12'h322, 12'h655, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h998, 12'h899, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h788, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h887, 12'h878, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h899, 12'h989, 12'h899, 12'h999, 12'h988, 12'h999, 12'h899, 12'h998, 12'h898, 12'h999, 12'h999, 12'h989, 12'h999, 12'h999, 12'h777, 12'h667, 12'h666, 12'hAAA, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFEE, 12'hDCC, 12'hCBA, 12'hCAA, 12'hDA9, 12'hEAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD98, 12'hC98, 12'hC98, 12'hC98, 12'hB98, 12'hB88, 12'hB87, 12'hB88, 12'hB88, 12'hB88, 12'hA88, 12'hA88, 12'hA88, 12'h977, 12'h977, 12'hA77, 12'hA88, 12'h977, 12'h977, 12'h987, 12'hA78, 12'h977, 12'h977, 12'h977, 12'h977, 12'h977, 12'h966, 12'h976, 12'h966, 12'h966, 12'h967, 12'h866, 12'h866, 12'h755, 12'h655, 12'h534, 12'h533, 12'h433, 12'h423, 12'h422, 12'h322, 12'h323, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h333, 12'h988, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h899, 12'h989, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h777, 12'h887, 12'h888, 12'h787, 12'h878, 12'h888, 12'h888, 12'h877, 12'h888, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h998, 12'h889, 12'h999, 12'h999, 12'h998, 12'h999, 12'h898, 12'h989, 12'h998, 12'h888, 12'h888, 12'h988, 12'h999, 12'h889, 12'h999, 12'h999, 12'h778, 12'h666, 12'h767, 12'h555, 12'h9AA, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFEE, 12'hDBB, 12'hCAA, 12'hDAA, 12'hDAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hC98, 12'hC98, 12'hD98, 12'hC98, 12'hC98, 12'hB87, 12'hB87, 12'hB87, 12'hA87, 12'hB88, 12'hB98, 12'hA98, 12'hA88, 12'hA88, 12'h988, 12'h987, 12'h977, 12'h977, 12'h866, 12'h866, 12'h866, 12'h866, 12'h755, 12'h755, 12'h755, 12'h755, 12'h755, 12'h745, 12'h644, 12'h644, 12'h644, 12'h644, 12'h544, 12'h533, 12'h433, 12'h423, 12'h322, 12'h323, 12'h432, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h322, 12'h322, 12'h333, 12'h333, 12'h322, 12'h544, 12'hAAA, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h777, 12'h878, 12'h888, 12'h787, 12'h878, 12'h787, 12'h888, 12'h788, 12'h878, 12'h887, 12'h888, 12'h778, 12'h787, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h999, 12'h888, 12'h899, 12'h988, 12'h999, 12'h999, 12'h999, 12'h999, 12'h989, 12'h898, 12'h999, 12'h998, 12'h888, 12'h998, 12'h888, 12'h999, 12'h999, 12'h888, 12'h667, 12'h666, 12'h556, 12'h667, 12'h678, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFDD, 12'hDBB, 12'hCAA, 12'hCAA, 12'hDAA, 12'hDA9, 12'hDA9, 12'hDA9, 12'hD99, 12'hD98, 12'hC88, 12'hC88, 12'hB88, 12'hB88, 12'hB87, 12'hA88, 12'hB88, 12'hB88, 12'hA88, 12'hA88, 12'hA88, 12'hA87, 12'hA87, 12'h977, 12'h977, 12'h977, 12'h877, 12'h866, 12'h766, 12'h755, 12'h655, 12'h645, 12'h645, 12'h644, 12'h544, 12'h534, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h323, 12'h322, 12'h322, 12'h323, 12'h322, 12'h322, 12'h332, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h333, 12'h322, 12'h322, 12'h776, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h9A9, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h787, 12'h878, 12'h888, 12'h888, 12'h877, 12'h787, 12'h878, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h999, 12'h889, 12'h888, 12'h998, 12'h999, 12'h888, 12'h998, 12'h999, 12'h899, 12'h998, 12'h989, 12'h899, 12'h998, 12'h899, 12'h898, 12'h989, 12'h888, 12'h777, 12'h667, 12'h556, 12'h556, 12'h656, 12'h667, 12'h556, 12'hCCD, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hDCB, 12'hB99, 12'hCAA, 12'hDBA, 12'hDA9, 12'hDA9, 12'hD99, 12'hD98, 12'hC98, 12'hB88, 12'hB87, 12'hB87, 12'hB88, 12'hB87, 12'hB87, 12'hA87, 12'hA87, 12'hA87, 12'hA87, 12'hA87, 12'h977, 12'h987, 12'h977, 12'h977, 12'h977, 12'h877, 12'h866, 12'h766, 12'h755, 12'h755, 12'h644, 12'h644, 12'h544, 12'h544, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h332, 12'h332, 12'h323, 12'h322, 12'h322, 12'h323, 12'h322, 12'h323, 12'h323, 12'h322, 12'h333, 12'h322, 12'h322, 12'h222, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h999, 12'h999, 12'hAA9, 12'hA99, 12'h9A9, 12'hAA9, 12'hAA9, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAA9, 12'h9A9, 12'h999, 12'h9A9, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h9A9,
		12'h888, 12'h777, 12'h787, 12'h888, 12'h878, 12'h788, 12'h877, 12'h777, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h898, 12'h999, 12'h999, 12'h999, 12'h888, 12'h998, 12'h999, 12'h899, 12'h989, 12'h999, 12'h998, 12'h998, 12'h889, 12'h999, 12'h988, 12'h888, 12'h998, 12'h888, 12'h666, 12'h566, 12'h656, 12'h556, 12'h556, 12'h557, 12'h667, 12'h445, 12'h456, 12'hDEE, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFDD, 12'hDBB, 12'hB99, 12'hC99, 12'hDA9, 12'hD99, 12'hD99, 12'hC99, 12'hC98, 12'hC88, 12'hC88, 12'hB87, 12'hB87, 12'hB77, 12'hB77, 12'hB77, 12'hA77, 12'hA77, 12'h977, 12'h977, 12'h976, 12'h976, 12'h976, 12'h977, 12'h966, 12'h866, 12'h866, 12'h755, 12'h755, 12'h655, 12'h644, 12'h644, 12'h544, 12'h534, 12'h533, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h332, 12'h322, 12'h323, 12'h322, 12'h322, 12'h322, 12'h423, 12'h322, 12'h433, 12'h322, 12'h332, 12'h344, 12'h999, 12'h9A9, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hA99, 12'hAAA, 12'h999, 12'hAA9, 12'hAA9, 12'h9A9, 12'h9A9, 12'h999, 12'h9A9, 12'h9A9,
		12'h888, 12'h878, 12'h888, 12'h888, 12'h778, 12'h888, 12'h888, 12'h778, 12'h888, 12'h877, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h999, 12'h888, 12'h999, 12'h999, 12'h888, 12'h989, 12'h999, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h888, 12'h999, 12'h889, 12'h888, 12'h667, 12'h656, 12'h667, 12'h657, 12'h556, 12'h556, 12'h556, 12'h556, 12'h555, 12'h556, 12'h456, 12'hCDE, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEDD, 12'hDAB, 12'hB99, 12'hC99, 12'hDA9, 12'hD99, 12'hD98, 12'hC88, 12'hB87, 12'hB76, 12'hB77, 12'hB87, 12'hB87, 12'hB87, 12'hB88, 12'hA87, 12'hA77, 12'hA77, 12'h976, 12'h976, 12'h966, 12'h866, 12'h866, 12'h866, 12'h755, 12'h755, 12'h644, 12'h644, 12'h544, 12'h543, 12'h533, 12'h533, 12'h433, 12'h433, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h422, 12'h322, 12'h322, 12'h433, 12'h323, 12'h222, 12'h777, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'hAA9, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h9A9, 12'h999, 12'h9A9, 12'h999, 12'hAAA, 12'h99A, 12'hA9A, 12'hAA9, 12'h9A9, 12'hAAA, 12'h999, 12'h9A9,
		12'h888, 12'h888, 12'h877, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h989, 12'h898, 12'h989, 12'h999, 12'h999, 12'h898, 12'h889, 12'h998, 12'h998, 12'h889, 12'h998, 12'h999, 12'h888, 12'h889, 12'h999, 12'h888, 12'h777, 12'h777, 12'h667, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h445, 12'h545, 12'h445, 12'h555, 12'h445, 12'h445, 12'hDFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFEF, 12'hFEE, 12'hDCC, 12'hC9A, 12'hC99, 12'hC98, 12'hD98, 12'hC98, 12'hC87, 12'hB87, 12'hB87, 12'hB87, 12'hB87, 12'hB88, 12'hB88, 12'hB87, 12'hA77, 12'hA77, 12'hA77, 12'h976, 12'h966, 12'h866, 12'h865, 12'h855, 12'h755, 12'h754, 12'h644, 12'h644, 12'h543, 12'h533, 12'h533, 12'h433, 12'h433, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h433, 12'h322, 12'h322, 12'h322, 12'h323, 12'h333, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'hA99, 12'h9A9, 12'hAA9, 12'h999, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'hAA9, 12'h999, 12'hAA9, 12'h9A9, 12'h99A, 12'hAA9, 12'h999, 12'h9A9, 12'hAA9, 12'h999, 12'h9A9, 12'h9A9, 12'h9A9, 12'h9A9, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h9A9, 12'h999, 12'h99A, 12'h999, 12'h999, 12'h9A9, 12'h999,
		12'h888, 12'h888, 12'h778, 12'h887, 12'h888, 12'h878, 12'h877, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h898, 12'h998, 12'h999, 12'h999, 12'h998, 12'h998, 12'h999, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h989, 12'h888, 12'h777, 12'h667, 12'h666, 12'h556, 12'h556, 12'h556, 12'h556, 12'h545, 12'h445, 12'h445, 12'h555, 12'h445, 12'h556, 12'h444, 12'h556, 12'h778, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hFFF, 12'hFEE, 12'hDBB, 12'hCAA, 12'hB98, 12'hC99, 12'hC98, 12'hC88, 12'hC87, 12'hC87, 12'hB77, 12'hB87, 12'hB88, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hA77, 12'hA77, 12'h976, 12'h966, 12'h966, 12'h865, 12'h855, 12'h855, 12'h754, 12'h644, 12'h644, 12'h543, 12'h533, 12'h433, 12'h422, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h433, 12'h423, 12'h433, 12'h433, 12'h322, 12'h322, 12'h444, 12'h888, 12'h9A9, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h9AA, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'h999, 12'hA99, 12'hA99, 12'hAA9, 12'h9A9, 12'hA99, 12'h9A9, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'hAAA, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h999,
		12'h888, 12'h878, 12'h888, 12'h788, 12'h878, 12'h788, 12'h888, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h998, 12'h998, 12'h899, 12'h998, 12'h999, 12'h999, 12'h988, 12'h998, 12'h999, 12'h998, 12'h998, 12'h999, 12'h889, 12'h888, 12'h777, 12'h666, 12'h666, 12'h667, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h445, 12'h445, 12'h546, 12'h434, 12'h556, 12'h334, 12'h445, 12'h445, 12'h445, 12'h9AB, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEE, 12'hFEF, 12'hDCC, 12'hC99, 12'hC99, 12'hC99, 12'hC88, 12'hC98, 12'hC88, 12'hC88, 12'hB87, 12'hC88, 12'hC88, 12'hC88, 12'hB88, 12'hB87, 12'hB77, 12'hA77, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h966, 12'h866, 12'h855, 12'h755, 12'h754, 12'h644, 12'h644, 12'h533, 12'h433, 12'h433, 12'h423, 12'h433, 12'h333, 12'h422, 12'h422, 12'h333, 12'h422, 12'h433, 12'h322, 12'h322, 12'h434, 12'h766, 12'h999, 12'h9AA, 12'hA99, 12'hAA9, 12'h9AA, 12'hA99, 12'h999, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'h99A, 12'hAA9, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAAA, 12'hAAA, 12'h99A, 12'hAA9, 12'hAA9, 12'h999, 12'h9A9, 12'h999, 12'hAA9, 12'h9A9, 12'h99A, 12'hAA9, 12'h9AA, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h887, 12'h877, 12'h888, 12'h888, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h998, 12'h999, 12'h888, 12'h999, 12'h999, 12'h888, 12'h999, 12'h999, 12'h777, 12'h667, 12'h666, 12'h666, 12'h556, 12'h556, 12'h555, 12'h556, 12'h556, 12'h555, 12'h545, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h345, 12'h689, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hFEF, 12'hEDD, 12'hCBA, 12'hB99, 12'hB88, 12'hC99, 12'hC98, 12'hB87, 12'hB77, 12'hB88, 12'hC88, 12'hC88, 12'hC88, 12'hC88, 12'hB87, 12'hB77, 12'hA76, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h966, 12'h966, 12'h855, 12'h755, 12'h745, 12'h644, 12'h644, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h322, 12'h422, 12'h433, 12'h433, 12'h323, 12'h554, 12'h666, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9AA, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'hAA9, 12'hAA9, 12'h999, 12'hAAA, 12'hAA9, 12'h9AA, 12'hAAA, 12'hAAA, 12'h9AA, 12'hA99, 12'h9AA, 12'hAA9, 12'hA9A, 12'h9A9, 12'h9A9, 12'hAAA, 12'h999, 12'h9AA, 12'h99A, 12'hA99, 12'h9A9, 12'h99A, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'h999, 12'h99A, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h788, 12'h878, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h988, 12'h988, 12'h898, 12'h988, 12'h998, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h989, 12'h888, 12'h777, 12'h666, 12'h667, 12'h657, 12'h556, 12'h556, 12'h556, 12'h555, 12'h545, 12'h545, 12'h545, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h435, 12'h334, 12'h345, 12'h345, 12'h335, 12'h457, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hEFF, 12'hFFF, 12'hEED, 12'hCBB, 12'hB99, 12'hB99, 12'hB98, 12'hB88, 12'hB77, 12'hB77, 12'hB88, 12'hB87, 12'hB87, 12'hC87, 12'hB88, 12'hB77, 12'hA77, 12'hA76, 12'hA76, 12'hA76, 12'hA66, 12'h966, 12'h966, 12'h855, 12'h855, 12'h755, 12'h644, 12'h634, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h322, 12'h423, 12'h433, 12'h323, 12'h433, 12'h666, 12'h766, 12'hAAA, 12'hAAA, 12'h999, 12'h9AA, 12'hA9A, 12'h999, 12'hAA9, 12'hAAA, 12'h999, 12'hA99, 12'h9A9, 12'h99A, 12'hA99, 12'h9AA, 12'h99A, 12'hAA9, 12'h999, 12'h999, 12'hAA9, 12'hAAA, 12'h999, 12'h9A9, 12'hAAA, 12'h99A, 12'hAA9, 12'hAAA, 12'hAAA, 12'h999, 12'hAA9, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'hA9A, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h989, 12'h999, 12'h898, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99A, 12'h999, 12'h999, 12'h667, 12'h556, 12'h666, 12'h667, 12'h556, 12'h556, 12'h556, 12'h556, 12'h545, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h545, 12'h546, 12'h445, 12'h445, 12'h445, 12'h445, 12'h435, 12'h334, 12'h344, 12'h334, 12'h345, 12'h8AB, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEE, 12'hEEE, 12'hFEE, 12'hEDC, 12'hB99, 12'hA88, 12'hB99, 12'hC99, 12'hB78, 12'hB88, 12'hC88, 12'hB88, 12'hB77, 12'hB87, 12'hC88, 12'hB87, 12'hB77, 12'hB77, 12'hA77, 12'hA76, 12'h966, 12'h966, 12'h865, 12'h855, 12'h744, 12'h644, 12'h633, 12'h533, 12'h433, 12'h423, 12'h433, 12'h433, 12'h433, 12'h433, 12'h322, 12'h544, 12'h767, 12'h777, 12'h999, 12'h9AA, 12'hAA9, 12'hAAA, 12'hAA9, 12'h99A, 12'hAAA, 12'hAA9, 12'hAAA, 12'h9AA, 12'hA99, 12'h9A9, 12'hA9A, 12'h999, 12'h9A9, 12'hAAA, 12'h999, 12'hAAA, 12'h999, 12'h9A9, 12'hAAA, 12'hA99, 12'h9A9, 12'hA9A, 12'h9A9, 12'hAAA, 12'hA9A, 12'h9A9, 12'hA99, 12'hAAA, 12'h9A9, 12'hA99, 12'h99A, 12'h9A9, 12'hAA9, 12'h9AA, 12'h999, 12'hAA9, 12'h9AA, 12'h99A, 12'hAA9, 12'h9AA, 12'h999, 12'hAAA, 12'h999, 12'h9A9, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h989, 12'h989, 12'h898, 12'h989, 12'h989, 12'h999, 12'h999, 12'h999, 12'h899, 12'h777, 12'h656, 12'h445, 12'h445, 12'h445, 12'h455, 12'h556, 12'h556, 12'h546, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h435, 12'h334, 12'h334, 12'h334, 12'h444, 12'h334, 12'h334, 12'h245, 12'h79A, 12'hDFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEEF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEEF, 12'hDEE, 12'hEEE, 12'hEEE, 12'hDCC, 12'hCAA, 12'hB99, 12'hB89, 12'hB88, 12'hB78, 12'hB77, 12'hB88, 12'hC88, 12'hC88, 12'hC88, 12'hB87, 12'hB77, 12'hA76, 12'hA76, 12'h966, 12'h966, 12'h865, 12'h855, 12'h644, 12'h643, 12'h533, 12'h533, 12'h433, 12'h433, 12'h433, 12'h433, 12'h422, 12'h322, 12'h655, 12'h766, 12'h777, 12'h666, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA99, 12'hAAA, 12'hAAA, 12'h9A9, 12'hA9A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'hAA9, 12'hAAA, 12'h9AA, 12'hA99, 12'hAAA, 12'h9AA, 12'hA99, 12'hAAA, 12'h9A9, 12'hAAA, 12'h9A9, 12'hAAA, 12'h9AA, 12'h999, 12'hA9A, 12'h9A9, 12'h999, 12'hA99, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'hA9A, 12'h9A9, 12'hA99, 12'h99A, 12'h999, 12'h999,
		12'h887, 12'h887, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h999, 12'h999, 12'h888, 12'h778, 12'h778, 12'h677, 12'h667, 12'h556, 12'h555, 12'h444, 12'h334, 12'h344, 12'h434, 12'h444, 12'h445, 12'h445, 12'h445, 12'h445, 12'h444, 12'h444, 12'h334, 12'h334, 12'h434, 12'h444, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h445, 12'h334, 12'h445, 12'h445, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h346, 12'h357, 12'hDFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFEF, 12'hEEF, 12'hEFF, 12'hEFF, 12'hEEE, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDED, 12'hEDD, 12'hDCC, 12'hA99, 12'hA88, 12'hB99, 12'hB88, 12'hB77, 12'hB77, 12'hB88, 12'hB88, 12'hB87, 12'hB87, 12'hB77, 12'hA76, 12'hA66, 12'h966, 12'h754, 12'h644, 12'h644, 12'h533, 12'h533, 12'h433, 12'h533, 12'h533, 12'h433, 12'h322, 12'h766, 12'h888, 12'h878, 12'h777, 12'h667, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'h9A9, 12'hAA9, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAA9, 12'h9A9, 12'h999, 12'hAA9, 12'h9A9, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAA9, 12'h9AA, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h888, 12'h888, 12'h998, 12'h888, 12'h888, 12'h888, 12'h988, 12'h999, 12'h888, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h445, 12'h445, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h334, 12'h334, 12'h444, 12'h445, 12'h445, 12'h334, 12'h444, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h444, 12'h444, 12'h444, 12'h445, 12'h334, 12'h334, 12'h434, 12'h445, 12'h435, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h679, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEEF, 12'hFEF, 12'hEFF, 12'hEEE, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDEE, 12'hDDE, 12'hDDD, 12'hEDD, 12'hDCC, 12'hCAA, 12'hB88, 12'hB88, 12'hC88, 12'hB87, 12'hB88, 12'hB88, 12'hB77, 12'hA77, 12'hA66, 12'h965, 12'h855, 12'h643, 12'h533, 12'h533, 12'h533, 12'h543, 12'h433, 12'h534, 12'h433, 12'h433, 12'h766, 12'h988, 12'h878, 12'h877, 12'h777, 12'h777, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'hAA9, 12'h9A9, 12'h9A9, 12'hA99, 12'h9A9, 12'hAA9, 12'hAAA, 12'hA9A, 12'hAA9, 12'hAAA, 12'hAAA, 12'hA99, 12'hAAA, 12'hAA9, 12'hAAA, 12'hA99, 12'h9A9, 12'hAAA, 12'hA99, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'hAA9, 12'h9AA, 12'h9A9, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h998, 12'h888, 12'h888, 12'h998, 12'h999, 12'h999, 12'h888, 12'h667, 12'h666, 12'h667, 12'h556, 12'h445, 12'h555, 12'h445, 12'h445, 12'h334, 12'h444, 12'h334, 12'h223, 12'h223, 12'h333, 12'h334, 12'h334, 12'h444, 12'h445, 12'h434, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h324, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h234, 12'h89B, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEEF, 12'hEFF, 12'hEEF, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDDE, 12'hEEE, 12'hDDD, 12'hDCC, 12'hDCC, 12'hDBB, 12'hA88, 12'hA88, 12'hB88, 12'hB88, 12'hB88, 12'hB77, 12'hA77, 12'h966, 12'h855, 12'h744, 12'h634, 12'h644, 12'h644, 12'h644, 12'h544, 12'h544, 12'h433, 12'h433, 12'h777, 12'h988, 12'h999, 12'h878, 12'h878, 12'h777, 12'h777, 12'hAAB, 12'hAAB, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h999, 12'h999, 12'hAA9, 12'hAAA, 12'h9A9, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'h9AA, 12'hA99, 12'h9AA, 12'h9AA, 12'hA99, 12'h9AA, 12'h999, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'hAAA, 12'hAAA, 12'h999, 12'h999, 12'hA99, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999,
		12'h889, 12'h888, 12'h999, 12'h999, 12'h889, 12'h778, 12'h666, 12'h667, 12'h667, 12'h666, 12'h556, 12'h545, 12'h445, 12'h445, 12'h334, 12'h334, 12'h333, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h334, 12'h333, 12'h334, 12'h334, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h323, 12'h223, 12'h344, 12'h234, 12'h78A, 12'hDFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFEF, 12'hEFF, 12'hFFF, 12'hEEF, 12'hFFF, 12'hFFF, 12'hEEF, 12'hEEF, 12'hEEE, 12'hDEE, 12'hDEE, 12'hDDE, 12'hDDE, 12'hDDD, 12'hDCD, 12'hDCC, 12'hDCC, 12'hBAB, 12'hB99, 12'h977, 12'h966, 12'h977, 12'h966, 12'h855, 12'h744, 12'h744, 12'h643, 12'h644, 12'h644, 12'h645, 12'h545, 12'h433, 12'h656, 12'h988, 12'hA9A, 12'hA9A, 12'h999, 12'h888, 12'h888, 12'h777, 12'h777, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAA9, 12'h9A9, 12'hA99, 12'h999, 12'hAAA, 12'hA99, 12'h9AA, 12'hAA9, 12'hAA9, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'h9A9, 12'hA99, 12'hAAA, 12'h9A9, 12'hA99, 12'h9AA, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h999, 12'hAAA, 12'hAA9, 12'h999, 12'h99A, 12'h9A9, 12'hA99, 12'h99A, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h999, 12'h889, 12'h878, 12'h777, 12'h666, 12'h666, 12'h667, 12'h666, 12'h656, 12'h556, 12'h445, 12'h445, 12'h445, 12'h334, 12'h333, 12'h223, 12'h223, 12'h223, 12'h323, 12'h223, 12'h223, 12'h223, 12'h333, 12'h334, 12'h344, 12'h334, 12'h334, 12'h333, 12'h223, 12'h223, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h434, 12'h334, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h334, 12'h334, 12'h233, 12'h345, 12'h234, 12'h568, 12'hDFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFEF, 12'hFFF, 12'hEEF, 12'hEEF, 12'hEEF, 12'hEEF, 12'hDDE, 12'hDDE, 12'hDDD, 12'hCDD, 12'hCCD, 12'hCCC, 12'hCCC, 12'hDBC, 12'hB99, 12'h877, 12'h856, 12'h855, 12'h644, 12'h744, 12'h633, 12'h644, 12'h755, 12'h644, 12'h544, 12'h544, 12'h999, 12'hBAB, 12'hBAB, 12'hBBB, 12'h999, 12'h999, 12'h889, 12'h888, 12'h888, 12'h666, 12'hAAA, 12'h99A, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'hA99, 12'h999, 12'hAA9, 12'hA99, 12'h999, 12'hAAA, 12'hAAA, 12'h999, 12'h9A9, 12'hA9A, 12'hAA9, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hA99, 12'h999, 12'h999, 12'h999, 12'h999,
		12'h556, 12'h666, 12'h666, 12'h667, 12'h667, 12'h666, 12'h556, 12'h556, 12'h555, 12'h445, 12'h444, 12'h334, 12'h334, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h333, 12'h334, 12'h434, 12'h333, 12'h334, 12'h333, 12'h223, 12'h223, 12'h223, 12'h233, 12'h333, 12'h334, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h224, 12'h323, 12'h223, 12'h334, 12'h334, 12'h124, 12'h89B, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFEF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEEF, 12'hFFF, 12'hEEE, 12'hEEE, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDDE, 12'hDDE, 12'hDDD, 12'hCDD, 12'hCCC, 12'hCCC, 12'hCCC, 12'hCCC, 12'hBAA, 12'hA99, 12'h755, 12'h644, 12'h644, 12'h544, 12'h655, 12'h644, 12'h444, 12'h655, 12'hAAA, 12'hCCC, 12'hCCC, 12'hCCC, 12'hAAB, 12'hA9A, 12'h999, 12'h999, 12'h889, 12'h878, 12'h777, 12'h999, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'h9A9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'h9AA, 12'h9AA, 12'hA99, 12'h9A9, 12'h999, 12'hAA9, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h9AA, 12'hAA9, 12'h999, 12'hAAA, 12'hAA9, 12'h999, 12'h999,
		12'h667, 12'h667, 12'h667, 12'h556, 12'h546, 12'h545, 12'h445, 12'h445, 12'h444, 12'h334, 12'h334, 12'h333, 12'h323, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h122, 12'h223, 12'h223, 12'h223, 12'h333, 12'h334, 12'h344, 12'h334, 12'h334, 12'h223, 12'h233, 12'h223, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h223, 12'h223, 12'h233, 12'h223, 12'h334, 12'h345, 12'hABD, 12'hDFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEEF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFE, 12'hEEE, 12'hEEF, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDEE, 12'hDDE, 12'hCDD, 12'hCDD, 12'hCDD, 12'hCCD, 12'hCCC, 12'hCBC, 12'hBBB, 12'hAAA, 12'h766, 12'h433, 12'h655, 12'h544, 12'h766, 12'hA99, 12'hCBC, 12'hDDD, 12'hDDD, 12'hCCD, 12'hCCC, 12'hBBB, 12'hAAA, 12'h989, 12'h999, 12'h899, 12'h888, 12'h777, 12'h333, 12'h555, 12'h888, 12'h9AA, 12'hABA, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAA9, 12'hAA9, 12'hA9A, 12'hAAA, 12'hAA9, 12'hAAA, 12'h9AA, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'h9A9, 12'hA99, 12'h999, 12'h99A, 12'hAAA, 12'h9A9, 12'hAAA, 12'hA99, 12'h999,
		12'h556, 12'h546, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h223, 12'h333, 12'h334, 12'h334, 12'h334, 12'h333, 12'h223, 12'h223, 12'h223, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h324, 12'h334, 12'h334, 12'h223, 12'h333, 12'h223, 12'h333, 12'h223, 12'h345, 12'h99B, 12'hCDF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEEF, 12'hEEF, 12'hEEF, 12'hEEE, 12'hEEE, 12'hEEE, 12'hDDE, 12'hDDD, 12'hCDD, 12'hCDD, 12'hCCC, 12'hCCD, 12'hCCD, 12'hCCC, 12'hCBB, 12'h767, 12'h767, 12'h876, 12'h878, 12'hAAA, 12'h988, 12'h555, 12'h667, 12'hAAB, 12'hCCD, 12'hCCD, 12'hBAB, 12'hAAA, 12'h99A, 12'h999, 12'h888, 12'h888, 12'h777, 12'h222, 12'h222, 12'h111, 12'h111, 12'h444, 12'h999, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hABA, 12'hABA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9AA, 12'hAA9, 12'h9AA, 12'hAAA, 12'hA99, 12'hAAA, 12'h9A9, 12'hA9A, 12'hAAA, 12'h999, 12'h999, 12'h9A9, 12'hA9A, 12'h999, 12'h9AA, 12'hA99, 12'h999, 12'hAA9, 12'hA9A, 12'hAAA, 12'hAA9, 12'hA9A, 12'hAAA,
		12'h555, 12'h445, 12'h445, 12'h445, 12'h444, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h113, 12'h212, 12'h222, 12'h223, 12'h223, 12'h223, 12'h334, 12'h323, 12'h334, 12'h333, 12'h223, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h333, 12'h223, 12'h223, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h223, 12'h223, 12'h334, 12'h223, 12'h223, 12'h323, 12'h234, 12'h334, 12'h224, 12'h89B, 12'hCCF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFEF, 12'hEFF, 12'hFFF, 12'hEEF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hEEE, 12'hEEE, 12'hDEE, 12'hDDD, 12'hDDD, 12'hCDD, 12'hCDD, 12'hDDD, 12'hCCC, 12'hDDD, 12'h778, 12'h222, 12'h544, 12'h444, 12'h334, 12'h333, 12'h212, 12'h222, 12'h212, 12'h001, 12'h323, 12'h777, 12'hCCC, 12'hAAA, 12'hAAA, 12'h999, 12'h999, 12'h889, 12'h777, 12'h222, 12'h111, 12'h112, 12'h122, 12'h111, 12'h111, 12'h122, 12'h444, 12'h787, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'hAAA, 12'h9A9, 12'hAAA, 12'hAA9, 12'hAAA, 12'h9A9, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'h99A, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'hAA9, 12'h9AA, 12'hAA9, 12'hAAA, 12'h9AA, 12'hAA9, 12'hAAA, 12'h9A9, 12'hA99, 12'h999, 12'h999, 12'hA99, 12'hAAA, 12'hAAA,
		12'h445, 12'h445, 12'h444, 12'h334, 12'h334, 12'h334, 12'h333, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h222, 12'h123, 12'h222, 12'h213, 12'h122, 12'h222, 12'h223, 12'h223, 12'h334, 12'h334, 12'h334, 12'h333, 12'h233, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h333, 12'h323, 12'h233, 12'h223, 12'h223, 12'h324, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h223, 12'h223, 12'h223, 12'h223, 12'h323, 12'h223, 12'h223, 12'h334, 12'h334, 12'h334, 12'h234, 12'h99B, 12'hCDF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hEEF, 12'hEEE, 12'hDEE, 12'hDEE, 12'hDDE, 12'hDDD, 12'hDEE, 12'hCDD, 12'hDDD, 12'h999, 12'h111, 12'h111, 12'h222, 12'h222, 12'h111, 12'h212, 12'h112, 12'h112, 12'h111, 12'h222, 12'h112, 12'h111, 12'h223, 12'hAAB, 12'hBBC, 12'h99A, 12'h999, 12'h888, 12'h777, 12'h223, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h333, 12'h666, 12'h999, 12'hAAA, 12'hAAA, 12'h999, 12'h9A9, 12'h999, 12'h999, 12'h999, 12'h9A9, 12'h9A9, 12'hAAA, 12'h9A9, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAA9, 12'h9AA, 12'hAAA, 12'hAA9, 12'h999, 12'h9A9, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'hAA9, 12'h999, 12'hA9A, 12'h999, 12'hAAA, 12'hAAA, 12'h9A9, 12'h9AA, 12'hA9A, 12'h9A9, 12'hAA9,
		12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h233, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h233, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h223, 12'h223, 12'h323, 12'h333, 12'h334, 12'h334, 12'h333, 12'h223, 12'h323, 12'h323, 12'h323, 12'h323, 12'h334, 12'h334, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h445, 12'hBBC, 12'hBCE, 12'hDEF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hFFF, 12'hEFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hEEF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hEEF, 12'hEEE, 12'hDEE, 12'hDEE, 12'hDDD, 12'hCCC, 12'h333, 12'h111, 12'h222, 12'h112, 12'h111, 12'h212, 12'h222, 12'h222, 12'h222, 12'h323, 12'h222, 12'h223, 12'h222, 12'h111, 12'h222, 12'h111, 12'h434, 12'hAAA, 12'hAAA, 12'h888, 12'h777, 12'h223, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h212, 12'h222, 12'h112, 12'h112, 12'h111, 12'h222, 12'h444, 12'h555, 12'h999, 12'h999, 12'hAAA, 12'h999, 12'h999, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9AA, 12'h9AA, 12'h9AA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hA99, 12'h999, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h999, 12'h999, 12'hA99, 12'hA99, 12'hAA9, 12'hAA9, 12'h999, 12'h999,
		12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h333, 12'h334, 12'h334, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h323, 12'h323, 12'h333, 12'h223, 12'h223, 12'h323, 12'h323, 12'h334, 12'h334, 12'h334, 12'h334, 12'h223, 12'h333, 12'h233, 12'h233, 12'h344, 12'h89A, 12'hBCD, 12'hDEF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hFFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEFF, 12'hEEF, 12'hEEE, 12'hEEE, 12'hAAA, 12'h333, 12'h222, 12'h222, 12'h222, 12'h112, 12'h222, 12'h222, 12'h222, 12'h212, 12'h223, 12'h112, 12'h212, 12'h112, 12'h212, 12'h223, 12'h112, 12'h222, 12'h222, 12'h111, 12'h666, 12'hA9A, 12'h888, 12'h222, 12'h001, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h112, 12'h112, 12'h112, 12'h111, 12'h111, 12'h112, 12'h222, 12'h111, 12'h222, 12'h454, 12'h666, 12'h888, 12'hAAA, 12'hAA9, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'h9A9, 12'h9A9, 12'h999, 12'h999, 12'h9A9, 12'hAA9, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAAA, 12'hAA9, 12'hA99, 12'hA99, 12'hA99, 12'hA99, 12'h999, 12'h999, 12'h999,};

	assign rgb_colour = array[160*v_count_n+h_count_n];
endmodule